module crc32 ( gnd, vdd, data_in, crc_en, rst, clk, crc_out);

input gnd, vdd;
input crc_en;
input rst;
input clk;
input [7:0] data_in;
output [31:0] crc_out;

BUFX4 BUFX4_1 ( .A(_539__31_), .Y(_539__31_bF_buf3) );
BUFX4 BUFX4_2 ( .A(_539__31_), .Y(_539__31_bF_buf2) );
BUFX4 BUFX4_3 ( .A(_539__31_), .Y(_539__31_bF_buf1) );
BUFX4 BUFX4_4 ( .A(_539__31_), .Y(_539__31_bF_buf0) );
BUFX4 BUFX4_5 ( .A(_539__28_), .Y(_539__28_bF_buf3) );
BUFX4 BUFX4_6 ( .A(_539__28_), .Y(_539__28_bF_buf2) );
BUFX4 BUFX4_7 ( .A(_539__28_), .Y(_539__28_bF_buf1) );
BUFX4 BUFX4_8 ( .A(_539__28_), .Y(_539__28_bF_buf0) );
BUFX2 BUFX2_1 ( .A(clk), .Y(clk_bF_buf4) );
BUFX2 BUFX2_2 ( .A(clk), .Y(clk_bF_buf3) );
BUFX2 BUFX2_3 ( .A(clk), .Y(clk_bF_buf2) );
BUFX2 BUFX2_4 ( .A(clk), .Y(clk_bF_buf1) );
BUFX2 BUFX2_5 ( .A(clk), .Y(clk_bF_buf0) );
BUFX4 BUFX4_9 ( .A(crc_en), .Y(crc_en_bF_buf4) );
BUFX4 BUFX4_10 ( .A(crc_en), .Y(crc_en_bF_buf3) );
BUFX4 BUFX4_11 ( .A(crc_en), .Y(crc_en_bF_buf2) );
BUFX4 BUFX4_12 ( .A(crc_en), .Y(crc_en_bF_buf1) );
BUFX4 BUFX4_13 ( .A(crc_en), .Y(crc_en_bF_buf0) );
BUFX4 BUFX4_14 ( .A(_540_), .Y(_540__bF_buf4) );
BUFX4 BUFX4_15 ( .A(_540_), .Y(_540__bF_buf3) );
BUFX4 BUFX4_16 ( .A(_540_), .Y(_540__bF_buf2) );
BUFX4 BUFX4_17 ( .A(_540_), .Y(_540__bF_buf1) );
BUFX4 BUFX4_18 ( .A(_540_), .Y(_540__bF_buf0) );
BUFX4 BUFX4_19 ( .A(_539__30_), .Y(_539__30_bF_buf3) );
BUFX4 BUFX4_20 ( .A(_539__30_), .Y(_539__30_bF_buf2) );
BUFX4 BUFX4_21 ( .A(_539__30_), .Y(_539__30_bF_buf1) );
BUFX4 BUFX4_22 ( .A(_539__30_), .Y(_539__30_bF_buf0) );
BUFX4 BUFX4_23 ( .A(data_in[3]), .Y(data_in_3_bF_buf3) );
BUFX4 BUFX4_24 ( .A(data_in[3]), .Y(data_in_3_bF_buf2) );
BUFX4 BUFX4_25 ( .A(data_in[3]), .Y(data_in_3_bF_buf1) );
BUFX4 BUFX4_26 ( .A(data_in[3]), .Y(data_in_3_bF_buf0) );
BUFX4 BUFX4_27 ( .A(_516_), .Y(_516__bF_buf5) );
BUFX4 BUFX4_28 ( .A(_516_), .Y(_516__bF_buf4) );
BUFX4 BUFX4_29 ( .A(_516_), .Y(_516__bF_buf3) );
BUFX4 BUFX4_30 ( .A(_516_), .Y(_516__bF_buf2) );
BUFX4 BUFX4_31 ( .A(_516_), .Y(_516__bF_buf1) );
BUFX4 BUFX4_32 ( .A(_516_), .Y(_516__bF_buf0) );
BUFX4 BUFX4_33 ( .A(_539__29_), .Y(_539__29_bF_buf3) );
BUFX4 BUFX4_34 ( .A(_539__29_), .Y(_539__29_bF_buf2) );
BUFX4 BUFX4_35 ( .A(_539__29_), .Y(_539__29_bF_buf1) );
BUFX4 BUFX4_36 ( .A(_539__29_), .Y(_539__29_bF_buf0) );
AOI22X1 AOI22X1_1 ( .A(_524_), .B(_527_), .C(_533_), .D(_536_), .Y(_537_) );
NAND2X1 NAND2X1_1 ( .A(_524_), .B(_527_), .Y(_538_) );
NAND2X1 NAND2X1_2 ( .A(_539__31_bF_buf3), .B(_535_), .Y(_1_) );
NAND2X1 NAND2X1_3 ( .A(_534_), .B(_532_), .Y(_2_) );
AOI21X1 AOI21X1_1 ( .A(_1_), .B(_2_), .C(_538_), .Y(_3_) );
NAND2X1 NAND2X1_4 ( .A(data_in[6]), .B(data_in[7]), .Y(_4_) );
INVX2 INVX2_1 ( .A(data_in[6]), .Y(_5_) );
INVX2 INVX2_2 ( .A(data_in[7]), .Y(_6_) );
NAND2X1 NAND2X1_5 ( .A(_5_), .B(_6_), .Y(_7_) );
NAND2X1 NAND2X1_6 ( .A(_4_), .B(_7_), .Y(_8_) );
OAI21X1 OAI21X1_1 ( .A(_537_), .B(_3_), .C(_8_), .Y(_9_) );
NAND3X1 NAND3X1_1 ( .A(_1_), .B(_2_), .C(_538_), .Y(_10_) );
XOR2X1 XOR2X1_1 ( .A(_539__30_bF_buf3), .B(data_in[1]), .Y(_11_) );
NAND2X1 NAND2X1_7 ( .A(_539__24_), .B(_11_), .Y(_12_) );
INVX2 INVX2_3 ( .A(_539__24_), .Y(_13_) );
XNOR2X1 XNOR2X1_1 ( .A(_539__30_bF_buf2), .B(data_in[1]), .Y(_14_) );
NAND2X1 NAND2X1_8 ( .A(_13_), .B(_14_), .Y(_15_) );
NAND2X1 NAND2X1_9 ( .A(_15_), .B(_12_), .Y(_16_) );
NAND3X1 NAND3X1_2 ( .A(_533_), .B(_536_), .C(_16_), .Y(_17_) );
XOR2X1 XOR2X1_2 ( .A(data_in[6]), .B(data_in[7]), .Y(_18_) );
NAND3X1 NAND3X1_3 ( .A(_18_), .B(_10_), .C(_17_), .Y(_19_) );
NAND3X1 NAND3X1_4 ( .A(crc_en_bF_buf4), .B(_19_), .C(_9_), .Y(_20_) );
OAI21X1 OAI21X1_2 ( .A(crc_en_bF_buf3), .B(_521_), .C(_20_), .Y(_0__1_) );
INVX1 INVX1_1 ( .A(_539__2_), .Y(_21_) );
XNOR2X1 XNOR2X1_2 ( .A(_539__26_), .B(data_in[2]), .Y(_22_) );
XNOR2X1 XNOR2X1_3 ( .A(_18_), .B(_22_), .Y(_23_) );
NAND3X1 NAND3X1_5 ( .A(_23_), .B(_10_), .C(_17_), .Y(_24_) );
XNOR2X1 XNOR2X1_4 ( .A(_8_), .B(_22_), .Y(_25_) );
OAI21X1 OAI21X1_3 ( .A(_537_), .B(_3_), .C(_25_), .Y(_26_) );
NAND3X1 NAND3X1_6 ( .A(crc_en_bF_buf2), .B(_24_), .C(_26_), .Y(_27_) );
OAI21X1 OAI21X1_4 ( .A(crc_en_bF_buf1), .B(_21_), .C(_27_), .Y(_0__2_) );
NAND2X1 NAND2X1_10 ( .A(_539__3_), .B(_516__bF_buf5), .Y(_28_) );
INVX2 INVX2_4 ( .A(_539__26_), .Y(_29_) );
NAND2X1 NAND2X1_11 ( .A(_539__25_), .B(_29_), .Y(_30_) );
NAND2X1 NAND2X1_12 ( .A(_539__26_), .B(_530_), .Y(_31_) );
NAND2X1 NAND2X1_13 ( .A(_30_), .B(_31_), .Y(_32_) );
XNOR2X1 XNOR2X1_5 ( .A(data_in[2]), .B(data_in_3_bF_buf3), .Y(_33_) );
NAND2X1 NAND2X1_14 ( .A(_33_), .B(_32_), .Y(_34_) );
NAND2X1 NAND2X1_15 ( .A(_530_), .B(_29_), .Y(_35_) );
NAND2X1 NAND2X1_16 ( .A(_539__25_), .B(_539__26_), .Y(_36_) );
NAND2X1 NAND2X1_17 ( .A(_36_), .B(_35_), .Y(_37_) );
XOR2X1 XOR2X1_3 ( .A(data_in[2]), .B(data_in_3_bF_buf2), .Y(_38_) );
NAND2X1 NAND2X1_18 ( .A(_38_), .B(_37_), .Y(_39_) );
NOR2X1 NOR2X1_1 ( .A(data_in[1]), .B(_539__27_), .Y(_40_) );
NAND2X1 NAND2X1_19 ( .A(data_in[1]), .B(_539__27_), .Y(_41_) );
INVX1 INVX1_2 ( .A(_41_), .Y(_42_) );
OAI21X1 OAI21X1_5 ( .A(_40_), .B(_42_), .C(_539__31_bF_buf2), .Y(_43_) );
INVX1 INVX1_3 ( .A(_40_), .Y(_44_) );
NAND3X1 NAND3X1_7 ( .A(_534_), .B(_41_), .C(_44_), .Y(_45_) );
AND2X2 AND2X2_1 ( .A(_45_), .B(_43_), .Y(_46_) );
NAND3X1 NAND3X1_8 ( .A(_34_), .B(_39_), .C(_46_), .Y(_47_) );
NOR2X1 NOR2X1_2 ( .A(_38_), .B(_37_), .Y(_48_) );
INVX1 INVX1_4 ( .A(_39_), .Y(_49_) );
NAND2X1 NAND2X1_20 ( .A(_43_), .B(_45_), .Y(_50_) );
OAI21X1 OAI21X1_6 ( .A(_48_), .B(_49_), .C(_50_), .Y(_51_) );
NAND3X1 NAND3X1_9 ( .A(data_in[7]), .B(_47_), .C(_51_), .Y(_52_) );
NAND3X1 NAND3X1_10 ( .A(_34_), .B(_39_), .C(_50_), .Y(_53_) );
OAI21X1 OAI21X1_7 ( .A(_48_), .B(_49_), .C(_46_), .Y(_54_) );
NAND3X1 NAND3X1_11 ( .A(_6_), .B(_53_), .C(_54_), .Y(_55_) );
NAND3X1 NAND3X1_12 ( .A(crc_en_bF_buf0), .B(_55_), .C(_52_), .Y(_56_) );
NAND2X1 NAND2X1_21 ( .A(_28_), .B(_56_), .Y(_0__3_) );
INVX1 INVX1_5 ( .A(_539__4_), .Y(_57_) );
XNOR2X1 XNOR2X1_6 ( .A(_539__30_bF_buf1), .B(data_in[0]), .Y(_58_) );
INVX2 INVX2_5 ( .A(data_in[2]), .Y(_59_) );
INVX2 INVX2_6 ( .A(_539__28_bF_buf3), .Y(_60_) );
NAND2X1 NAND2X1_22 ( .A(_59_), .B(_60_), .Y(_61_) );
NAND2X1 NAND2X1_23 ( .A(data_in[2]), .B(_539__28_bF_buf2), .Y(_62_) );
NAND2X1 NAND2X1_24 ( .A(_62_), .B(_61_), .Y(_63_) );
XOR2X1 XOR2X1_4 ( .A(_63_), .B(_58_), .Y(_64_) );
NOR2X1 NOR2X1_3 ( .A(_539__26_), .B(_13_), .Y(_65_) );
NOR2X1 NOR2X1_4 ( .A(_539__24_), .B(_29_), .Y(_66_) );
OAI21X1 OAI21X1_8 ( .A(_65_), .B(_66_), .C(_539__27_), .Y(_67_) );
INVX2 INVX2_7 ( .A(_539__27_), .Y(_68_) );
NOR2X1 NOR2X1_5 ( .A(_539__24_), .B(_539__26_), .Y(_69_) );
NOR2X1 NOR2X1_6 ( .A(_13_), .B(_29_), .Y(_70_) );
OAI21X1 OAI21X1_9 ( .A(_69_), .B(_70_), .C(_68_), .Y(_71_) );
NAND2X1 NAND2X1_25 ( .A(_67_), .B(_71_), .Y(_72_) );
INVX4 INVX4_1 ( .A(data_in[4]), .Y(_73_) );
XOR2X1 XOR2X1_5 ( .A(data_in[6]), .B(data_in_3_bF_buf1), .Y(_74_) );
OR2X2 OR2X2_1 ( .A(_74_), .B(_73_), .Y(_75_) );
NAND2X1 NAND2X1_26 ( .A(_73_), .B(_74_), .Y(_76_) );
NAND3X1 NAND3X1_13 ( .A(_75_), .B(_76_), .C(_72_), .Y(_77_) );
OAI21X1 OAI21X1_10 ( .A(_65_), .B(_66_), .C(_68_), .Y(_78_) );
OAI21X1 OAI21X1_11 ( .A(_69_), .B(_70_), .C(_539__27_), .Y(_79_) );
NAND2X1 NAND2X1_27 ( .A(_78_), .B(_79_), .Y(_80_) );
NAND2X1 NAND2X1_28 ( .A(data_in[6]), .B(data_in[4]), .Y(_81_) );
NAND2X1 NAND2X1_29 ( .A(_5_), .B(_73_), .Y(_82_) );
AND2X2 AND2X2_2 ( .A(_82_), .B(_81_), .Y(_83_) );
NAND2X1 NAND2X1_30 ( .A(data_in_3_bF_buf0), .B(_83_), .Y(_84_) );
INVX1 INVX1_6 ( .A(data_in_3_bF_buf3), .Y(_85_) );
NAND2X1 NAND2X1_31 ( .A(_81_), .B(_82_), .Y(_86_) );
NAND2X1 NAND2X1_32 ( .A(_85_), .B(_86_), .Y(_87_) );
NAND3X1 NAND3X1_14 ( .A(_84_), .B(_87_), .C(_80_), .Y(_88_) );
NAND3X1 NAND3X1_15 ( .A(_64_), .B(_77_), .C(_88_), .Y(_89_) );
XNOR2X1 XNOR2X1_7 ( .A(_63_), .B(_58_), .Y(_90_) );
AOI21X1 AOI21X1_2 ( .A(_84_), .B(_87_), .C(_80_), .Y(_91_) );
AOI21X1 AOI21X1_3 ( .A(_75_), .B(_76_), .C(_72_), .Y(_92_) );
OAI21X1 OAI21X1_12 ( .A(_91_), .B(_92_), .C(_90_), .Y(_93_) );
NAND3X1 NAND3X1_16 ( .A(crc_en_bF_buf4), .B(_89_), .C(_93_), .Y(_94_) );
OAI21X1 OAI21X1_13 ( .A(crc_en_bF_buf3), .B(_57_), .C(_94_), .Y(_0__4_) );
NAND2X1 NAND2X1_33 ( .A(_539__5_), .B(_516__bF_buf4), .Y(_95_) );
NOR3X1 NOR3X1_1 ( .A(_530_), .B(_522_), .C(_523_), .Y(_96_) );
OR2X2 OR2X2_2 ( .A(_539__30_bF_buf0), .B(_539__24_), .Y(_97_) );
NAND2X1 NAND2X1_34 ( .A(_539__30_bF_buf3), .B(_539__24_), .Y(_98_) );
AOI21X1 AOI21X1_4 ( .A(_97_), .B(_98_), .C(_539__25_), .Y(_99_) );
NAND2X1 NAND2X1_35 ( .A(_539__27_), .B(_60_), .Y(_100_) );
NAND2X1 NAND2X1_36 ( .A(_539__28_bF_buf1), .B(_68_), .Y(_101_) );
INVX1 INVX1_7 ( .A(_539__29_bF_buf3), .Y(_102_) );
NAND2X1 NAND2X1_37 ( .A(_539__31_bF_buf1), .B(_102_), .Y(_103_) );
NAND2X1 NAND2X1_38 ( .A(_539__29_bF_buf2), .B(_534_), .Y(_104_) );
AOI22X1 AOI22X1_2 ( .A(_100_), .B(_101_), .C(_103_), .D(_104_), .Y(_105_) );
NAND2X1 NAND2X1_39 ( .A(_539__27_), .B(_539__28_bF_buf0), .Y(_106_) );
BUFX2 BUFX2_6 ( .A(_539__0_), .Y(crc_out[0]) );
BUFX2 BUFX2_7 ( .A(_539__1_), .Y(crc_out[1]) );
BUFX2 BUFX2_8 ( .A(_539__2_), .Y(crc_out[2]) );
BUFX2 BUFX2_9 ( .A(_539__3_), .Y(crc_out[3]) );
BUFX2 BUFX2_10 ( .A(_539__4_), .Y(crc_out[4]) );
BUFX2 BUFX2_11 ( .A(_539__5_), .Y(crc_out[5]) );
BUFX2 BUFX2_12 ( .A(_539__6_), .Y(crc_out[6]) );
BUFX2 BUFX2_13 ( .A(_539__7_), .Y(crc_out[7]) );
BUFX2 BUFX2_14 ( .A(_539__8_), .Y(crc_out[8]) );
BUFX2 BUFX2_15 ( .A(_539__9_), .Y(crc_out[9]) );
BUFX2 BUFX2_16 ( .A(_539__10_), .Y(crc_out[10]) );
BUFX2 BUFX2_17 ( .A(_539__11_), .Y(crc_out[11]) );
BUFX2 BUFX2_18 ( .A(_539__12_), .Y(crc_out[12]) );
BUFX2 BUFX2_19 ( .A(_539__13_), .Y(crc_out[13]) );
BUFX2 BUFX2_20 ( .A(_539__14_), .Y(crc_out[14]) );
BUFX2 BUFX2_21 ( .A(_539__15_), .Y(crc_out[15]) );
BUFX2 BUFX2_22 ( .A(_539__16_), .Y(crc_out[16]) );
BUFX2 BUFX2_23 ( .A(_539__17_), .Y(crc_out[17]) );
BUFX2 BUFX2_24 ( .A(_539__18_), .Y(crc_out[18]) );
BUFX2 BUFX2_25 ( .A(_539__19_), .Y(crc_out[19]) );
BUFX2 BUFX2_26 ( .A(_539__20_), .Y(crc_out[20]) );
BUFX2 BUFX2_27 ( .A(_539__21_), .Y(crc_out[21]) );
BUFX2 BUFX2_28 ( .A(_539__22_), .Y(crc_out[22]) );
BUFX2 BUFX2_29 ( .A(_539__23_), .Y(crc_out[23]) );
BUFX2 BUFX2_30 ( .A(_539__24_), .Y(crc_out[24]) );
BUFX2 BUFX2_31 ( .A(_539__25_), .Y(crc_out[25]) );
BUFX2 BUFX2_32 ( .A(_539__26_), .Y(crc_out[26]) );
BUFX2 BUFX2_33 ( .A(_539__27_), .Y(crc_out[27]) );
BUFX2 BUFX2_34 ( .A(_539__28_bF_buf3), .Y(crc_out[28]) );
BUFX2 BUFX2_35 ( .A(_539__29_bF_buf1), .Y(crc_out[29]) );
BUFX2 BUFX2_36 ( .A(_539__30_bF_buf2), .Y(crc_out[30]) );
BUFX2 BUFX2_37 ( .A(_539__31_bF_buf0), .Y(crc_out[31]) );
DFFSR DFFSR_1 ( .CLK(clk_bF_buf4), .D(_0__0_), .Q(_539__0_), .R(vdd), .S(_540__bF_buf4) );
DFFSR DFFSR_2 ( .CLK(clk_bF_buf3), .D(_0__1_), .Q(_539__1_), .R(vdd), .S(_540__bF_buf3) );
DFFSR DFFSR_3 ( .CLK(clk_bF_buf2), .D(_0__2_), .Q(_539__2_), .R(vdd), .S(_540__bF_buf2) );
DFFSR DFFSR_4 ( .CLK(clk_bF_buf1), .D(_0__3_), .Q(_539__3_), .R(vdd), .S(_540__bF_buf1) );
DFFSR DFFSR_5 ( .CLK(clk_bF_buf0), .D(_0__4_), .Q(_539__4_), .R(vdd), .S(_540__bF_buf0) );
DFFSR DFFSR_6 ( .CLK(clk_bF_buf4), .D(_0__5_), .Q(_539__5_), .R(vdd), .S(_540__bF_buf4) );
DFFSR DFFSR_7 ( .CLK(clk_bF_buf3), .D(_0__6_), .Q(_539__6_), .R(vdd), .S(_540__bF_buf3) );
DFFSR DFFSR_8 ( .CLK(clk_bF_buf2), .D(_0__7_), .Q(_539__7_), .R(vdd), .S(_540__bF_buf2) );
DFFSR DFFSR_9 ( .CLK(clk_bF_buf1), .D(_0__8_), .Q(_539__8_), .R(vdd), .S(_540__bF_buf1) );
DFFSR DFFSR_10 ( .CLK(clk_bF_buf0), .D(_0__9_), .Q(_539__9_), .R(vdd), .S(_540__bF_buf0) );
DFFSR DFFSR_11 ( .CLK(clk_bF_buf4), .D(_0__10_), .Q(_539__10_), .R(vdd), .S(_540__bF_buf4) );
DFFSR DFFSR_12 ( .CLK(clk_bF_buf3), .D(_0__11_), .Q(_539__11_), .R(vdd), .S(_540__bF_buf3) );
DFFSR DFFSR_13 ( .CLK(clk_bF_buf2), .D(_0__12_), .Q(_539__12_), .R(vdd), .S(_540__bF_buf2) );
DFFSR DFFSR_14 ( .CLK(clk_bF_buf1), .D(_0__13_), .Q(_539__13_), .R(vdd), .S(_540__bF_buf1) );
DFFSR DFFSR_15 ( .CLK(clk_bF_buf0), .D(_0__14_), .Q(_539__14_), .R(vdd), .S(_540__bF_buf0) );
DFFSR DFFSR_16 ( .CLK(clk_bF_buf4), .D(_0__15_), .Q(_539__15_), .R(vdd), .S(_540__bF_buf4) );
DFFSR DFFSR_17 ( .CLK(clk_bF_buf3), .D(_0__16_), .Q(_539__16_), .R(vdd), .S(_540__bF_buf3) );
DFFSR DFFSR_18 ( .CLK(clk_bF_buf2), .D(_0__17_), .Q(_539__17_), .R(vdd), .S(_540__bF_buf2) );
DFFSR DFFSR_19 ( .CLK(clk_bF_buf1), .D(_0__18_), .Q(_539__18_), .R(vdd), .S(_540__bF_buf1) );
DFFSR DFFSR_20 ( .CLK(clk_bF_buf0), .D(_0__19_), .Q(_539__19_), .R(vdd), .S(_540__bF_buf0) );
DFFSR DFFSR_21 ( .CLK(clk_bF_buf4), .D(_0__20_), .Q(_539__20_), .R(vdd), .S(_540__bF_buf4) );
DFFSR DFFSR_22 ( .CLK(clk_bF_buf3), .D(_0__21_), .Q(_539__21_), .R(vdd), .S(_540__bF_buf3) );
DFFSR DFFSR_23 ( .CLK(clk_bF_buf2), .D(_0__22_), .Q(_539__22_), .R(vdd), .S(_540__bF_buf2) );
DFFSR DFFSR_24 ( .CLK(clk_bF_buf1), .D(_0__23_), .Q(_539__23_), .R(vdd), .S(_540__bF_buf1) );
DFFSR DFFSR_25 ( .CLK(clk_bF_buf0), .D(_0__24_), .Q(_539__24_), .R(vdd), .S(_540__bF_buf0) );
DFFSR DFFSR_26 ( .CLK(clk_bF_buf4), .D(_0__25_), .Q(_539__25_), .R(vdd), .S(_540__bF_buf4) );
DFFSR DFFSR_27 ( .CLK(clk_bF_buf3), .D(_0__26_), .Q(_539__26_), .R(vdd), .S(_540__bF_buf3) );
DFFSR DFFSR_28 ( .CLK(clk_bF_buf2), .D(_0__27_), .Q(_539__27_), .R(vdd), .S(_540__bF_buf2) );
DFFSR DFFSR_29 ( .CLK(clk_bF_buf1), .D(_0__28_), .Q(_539__28_), .R(vdd), .S(_540__bF_buf1) );
DFFSR DFFSR_30 ( .CLK(clk_bF_buf0), .D(_0__29_), .Q(_539__29_), .R(vdd), .S(_540__bF_buf0) );
DFFSR DFFSR_31 ( .CLK(clk_bF_buf4), .D(_0__30_), .Q(_539__30_), .R(vdd), .S(_540__bF_buf4) );
DFFSR DFFSR_32 ( .CLK(clk_bF_buf3), .D(_0__31_), .Q(_539__31_), .R(vdd), .S(_540__bF_buf3) );
OR2X2 OR2X2_3 ( .A(_539__27_), .B(_539__28_bF_buf2), .Y(_107_) );
NAND2X1 NAND2X1_40 ( .A(_539__31_bF_buf3), .B(_539__29_bF_buf0), .Y(_108_) );
OR2X2 OR2X2_4 ( .A(_539__31_bF_buf2), .B(_539__29_bF_buf3), .Y(_109_) );
AOI22X1 AOI22X1_3 ( .A(_107_), .B(_106_), .C(_108_), .D(_109_), .Y(_110_) );
OAI22X1 OAI22X1_1 ( .A(_96_), .B(_99_), .C(_110_), .D(_105_), .Y(_111_) );
AOI21X1 AOI21X1_5 ( .A(_97_), .B(_98_), .C(_530_), .Y(_112_) );
NOR3X1 NOR3X1_2 ( .A(_539__25_), .B(_522_), .C(_523_), .Y(_113_) );
AOI22X1 AOI22X1_4 ( .A(_109_), .B(_108_), .C(_100_), .D(_101_), .Y(_114_) );
AOI22X1 AOI22X1_5 ( .A(_107_), .B(_106_), .C(_103_), .D(_104_), .Y(_115_) );
OAI22X1 OAI22X1_2 ( .A(_112_), .B(_113_), .C(_114_), .D(_115_), .Y(_116_) );
AND2X2 AND2X2_3 ( .A(_111_), .B(_116_), .Y(_117_) );
NOR2X1 NOR2X1_7 ( .A(data_in[5]), .B(_5_), .Y(_118_) );
INVX4 INVX4_2 ( .A(data_in[5]), .Y(_119_) );
NOR2X1 NOR2X1_8 ( .A(data_in[6]), .B(_119_), .Y(_120_) );
NOR2X1 NOR2X1_9 ( .A(data_in[1]), .B(_529_), .Y(_121_) );
NOR2X1 NOR2X1_10 ( .A(data_in[0]), .B(_525_), .Y(_122_) );
OAI22X1 OAI22X1_3 ( .A(_118_), .B(_120_), .C(_121_), .D(_122_), .Y(_123_) );
AND2X2 AND2X2_4 ( .A(data_in[6]), .B(data_in[5]), .Y(_124_) );
NOR2X1 NOR2X1_11 ( .A(data_in[6]), .B(data_in[5]), .Y(_125_) );
AND2X2 AND2X2_5 ( .A(data_in[0]), .B(data_in[1]), .Y(_126_) );
NOR2X1 NOR2X1_12 ( .A(data_in[0]), .B(data_in[1]), .Y(_127_) );
OAI22X1 OAI22X1_4 ( .A(_125_), .B(_124_), .C(_126_), .D(_127_), .Y(_128_) );
NOR2X1 NOR2X1_13 ( .A(data_in[4]), .B(_85_), .Y(_129_) );
NOR2X1 NOR2X1_14 ( .A(data_in_3_bF_buf2), .B(_73_), .Y(_130_) );
OAI21X1 OAI21X1_14 ( .A(_129_), .B(_130_), .C(_6_), .Y(_131_) );
AND2X2 AND2X2_6 ( .A(data_in_3_bF_buf1), .B(data_in[4]), .Y(_132_) );
NOR2X1 NOR2X1_15 ( .A(data_in_3_bF_buf0), .B(data_in[4]), .Y(_133_) );
OAI21X1 OAI21X1_15 ( .A(_133_), .B(_132_), .C(data_in[7]), .Y(_134_) );
NAND2X1 NAND2X1_41 ( .A(_134_), .B(_131_), .Y(_135_) );
NAND3X1 NAND3X1_17 ( .A(_123_), .B(_128_), .C(_135_), .Y(_136_) );
NAND2X1 NAND2X1_42 ( .A(_128_), .B(_123_), .Y(_137_) );
NAND3X1 NAND3X1_18 ( .A(_131_), .B(_134_), .C(_137_), .Y(_138_) );
NAND3X1 NAND3X1_19 ( .A(_136_), .B(_138_), .C(_117_), .Y(_139_) );
NAND2X1 NAND2X1_43 ( .A(_116_), .B(_111_), .Y(_140_) );
AOI21X1 AOI21X1_6 ( .A(_131_), .B(_134_), .C(_137_), .Y(_141_) );
AOI21X1 AOI21X1_7 ( .A(_123_), .B(_128_), .C(_135_), .Y(_142_) );
OAI21X1 OAI21X1_16 ( .A(_142_), .B(_141_), .C(_140_), .Y(_143_) );
NAND3X1 NAND3X1_20 ( .A(crc_en_bF_buf2), .B(_143_), .C(_139_), .Y(_144_) );
NAND2X1 NAND2X1_44 ( .A(_95_), .B(_144_), .Y(_0__5_) );
NAND2X1 NAND2X1_45 ( .A(_539__6_), .B(_516__bF_buf3), .Y(_145_) );
XNOR2X1 XNOR2X1_8 ( .A(data_in[2]), .B(data_in[4]), .Y(_146_) );
NAND2X1 NAND2X1_46 ( .A(_108_), .B(_109_), .Y(_147_) );
NAND2X1 NAND2X1_47 ( .A(_147_), .B(_32_), .Y(_148_) );
NAND2X1 NAND2X1_48 ( .A(_103_), .B(_104_), .Y(_149_) );
NAND2X1 NAND2X1_49 ( .A(_37_), .B(_149_), .Y(_150_) );
NAND3X1 NAND3X1_21 ( .A(_146_), .B(_148_), .C(_150_), .Y(_151_) );
XOR2X1 XOR2X1_6 ( .A(data_in[2]), .B(data_in[4]), .Y(_152_) );
AOI22X1 AOI22X1_6 ( .A(_109_), .B(_108_), .C(_30_), .D(_31_), .Y(_153_) );
AOI22X1 AOI22X1_7 ( .A(_103_), .B(_104_), .C(_35_), .D(_36_), .Y(_154_) );
OAI21X1 OAI21X1_17 ( .A(_153_), .B(_154_), .C(_152_), .Y(_155_) );
NAND2X1 NAND2X1_50 ( .A(_155_), .B(_151_), .Y(_156_) );
XOR2X1 XOR2X1_7 ( .A(_539__28_bF_buf1), .B(data_in[5]), .Y(_157_) );
NOR2X1 NOR2X1_16 ( .A(_14_), .B(_8_), .Y(_158_) );
AOI21X1 AOI21X1_8 ( .A(_4_), .B(_7_), .C(_11_), .Y(_159_) );
OAI21X1 OAI21X1_18 ( .A(_159_), .B(_158_), .C(_157_), .Y(_160_) );
INVX1 INVX1_8 ( .A(_157_), .Y(_161_) );
NAND2X1 NAND2X1_51 ( .A(_11_), .B(_18_), .Y(_162_) );
NAND2X1 NAND2X1_52 ( .A(_14_), .B(_8_), .Y(_163_) );
NAND3X1 NAND3X1_22 ( .A(_161_), .B(_162_), .C(_163_), .Y(_164_) );
NAND3X1 NAND3X1_23 ( .A(_160_), .B(_164_), .C(_156_), .Y(_165_) );
NAND2X1 NAND2X1_53 ( .A(data_in[2]), .B(data_in[4]), .Y(_166_) );
NAND2X1 NAND2X1_54 ( .A(_59_), .B(_73_), .Y(_167_) );
AOI22X1 AOI22X1_8 ( .A(_30_), .B(_31_), .C(_166_), .D(_167_), .Y(_168_) );
INVX1 INVX1_9 ( .A(_168_), .Y(_169_) );
NAND2X1 NAND2X1_55 ( .A(_152_), .B(_37_), .Y(_170_) );
AOI21X1 AOI21X1_9 ( .A(_169_), .B(_170_), .C(_149_), .Y(_171_) );
NOR2X1 NOR2X1_17 ( .A(_146_), .B(_32_), .Y(_172_) );
NOR3X1 NOR3X1_3 ( .A(_147_), .B(_168_), .C(_172_), .Y(_173_) );
AOI21X1 AOI21X1_10 ( .A(_163_), .B(_162_), .C(_161_), .Y(_174_) );
NOR3X1 NOR3X1_4 ( .A(_157_), .B(_159_), .C(_158_), .Y(_175_) );
OAI22X1 OAI22X1_5 ( .A(_171_), .B(_173_), .C(_174_), .D(_175_), .Y(_176_) );
NAND3X1 NAND3X1_24 ( .A(crc_en_bF_buf1), .B(_176_), .C(_165_), .Y(_177_) );
NAND2X1 NAND2X1_56 ( .A(_145_), .B(_177_), .Y(_0__6_) );
NAND2X1 NAND2X1_57 ( .A(_539__7_), .B(_516__bF_buf2), .Y(_178_) );
XNOR2X1 XNOR2X1_9 ( .A(data_in[2]), .B(_539__29_bF_buf2), .Y(_179_) );
XOR2X1 XOR2X1_8 ( .A(data_in[0]), .B(_539__31_bF_buf1), .Y(_180_) );
NAND2X1 NAND2X1_58 ( .A(_179_), .B(_180_), .Y(_181_) );
XOR2X1 XOR2X1_9 ( .A(data_in[2]), .B(_539__29_bF_buf1), .Y(_182_) );
XNOR2X1 XNOR2X1_10 ( .A(data_in[0]), .B(_539__31_bF_buf0), .Y(_183_) );
NAND2X1 NAND2X1_59 ( .A(_183_), .B(_182_), .Y(_184_) );
XOR2X1 XOR2X1_10 ( .A(data_in_3_bF_buf3), .B(data_in[5]), .Y(_185_) );
AOI21X1 AOI21X1_11 ( .A(_181_), .B(_184_), .C(_185_), .Y(_186_) );
NAND2X1 NAND2X1_60 ( .A(_180_), .B(_182_), .Y(_187_) );
NAND2X1 NAND2X1_61 ( .A(_179_), .B(_183_), .Y(_188_) );
INVX1 INVX1_10 ( .A(_185_), .Y(_189_) );
AOI21X1 AOI21X1_12 ( .A(_187_), .B(_188_), .C(_189_), .Y(_190_) );
NAND3X1 NAND3X1_25 ( .A(_6_), .B(_67_), .C(_71_), .Y(_191_) );
NAND3X1 NAND3X1_26 ( .A(data_in[7]), .B(_78_), .C(_79_), .Y(_192_) );
NAND2X1 NAND2X1_62 ( .A(_191_), .B(_192_), .Y(_193_) );
OAI21X1 OAI21X1_19 ( .A(_186_), .B(_190_), .C(_193_), .Y(_194_) );
AOI21X1 AOI21X1_13 ( .A(_187_), .B(_188_), .C(_185_), .Y(_195_) );
AOI21X1 AOI21X1_14 ( .A(_184_), .B(_181_), .C(_189_), .Y(_196_) );
AND2X2 AND2X2_7 ( .A(_191_), .B(_192_), .Y(_197_) );
OAI21X1 OAI21X1_20 ( .A(_195_), .B(_196_), .C(_197_), .Y(_198_) );
NAND3X1 NAND3X1_27 ( .A(crc_en_bF_buf0), .B(_194_), .C(_198_), .Y(_199_) );
NAND2X1 NAND2X1_63 ( .A(_178_), .B(_199_), .Y(_0__7_) );
XNOR2X1 XNOR2X1_11 ( .A(data_in[0]), .B(_539__28_bF_buf0), .Y(_200_) );
NOR2X1 NOR2X1_18 ( .A(_539__25_), .B(_13_), .Y(_201_) );
NOR2X1 NOR2X1_19 ( .A(_539__24_), .B(_530_), .Y(_202_) );
OAI21X1 OAI21X1_21 ( .A(_201_), .B(_202_), .C(data_in[4]), .Y(_203_) );
NAND2X1 NAND2X1_64 ( .A(_13_), .B(_530_), .Y(_204_) );
NAND2X1 NAND2X1_65 ( .A(_539__24_), .B(_539__25_), .Y(_205_) );
NAND2X1 NAND2X1_66 ( .A(_205_), .B(_204_), .Y(_206_) );
NAND2X1 NAND2X1_67 ( .A(_73_), .B(_206_), .Y(_207_) );
NAND3X1 NAND3X1_28 ( .A(_200_), .B(_203_), .C(_207_), .Y(_208_) );
XOR2X1 XOR2X1_11 ( .A(data_in[0]), .B(_539__28_bF_buf3), .Y(_209_) );
NAND2X1 NAND2X1_68 ( .A(_203_), .B(_207_), .Y(_210_) );
NAND2X1 NAND2X1_69 ( .A(_209_), .B(_210_), .Y(_211_) );
NAND2X1 NAND2X1_70 ( .A(_41_), .B(_44_), .Y(_212_) );
XNOR2X1 XNOR2X1_12 ( .A(_539__0_), .B(data_in_3_bF_buf2), .Y(_213_) );
XNOR2X1 XNOR2X1_13 ( .A(_212_), .B(_213_), .Y(_214_) );
NAND3X1 NAND3X1_29 ( .A(_208_), .B(_214_), .C(_211_), .Y(_215_) );
OAI21X1 OAI21X1_22 ( .A(_201_), .B(_202_), .C(_200_), .Y(_216_) );
NAND2X1 NAND2X1_71 ( .A(_209_), .B(_206_), .Y(_217_) );
NAND3X1 NAND3X1_30 ( .A(_73_), .B(_216_), .C(_217_), .Y(_218_) );
NAND2X1 NAND2X1_72 ( .A(_216_), .B(_217_), .Y(_219_) );
NAND2X1 NAND2X1_73 ( .A(data_in[4]), .B(_219_), .Y(_220_) );
XOR2X1 XOR2X1_12 ( .A(_212_), .B(_213_), .Y(_221_) );
NAND3X1 NAND3X1_31 ( .A(_218_), .B(_221_), .C(_220_), .Y(_222_) );
NAND2X1 NAND2X1_74 ( .A(_215_), .B(_222_), .Y(_223_) );
NAND2X1 NAND2X1_75 ( .A(_539__8_), .B(_516__bF_buf1), .Y(_224_) );
OAI21X1 OAI21X1_23 ( .A(_516__bF_buf0), .B(_223_), .C(_224_), .Y(_0__8_) );
NAND2X1 NAND2X1_76 ( .A(_539__9_), .B(_516__bF_buf5), .Y(_225_) );
XOR2X1 XOR2X1_13 ( .A(_539__1_), .B(data_in[4]), .Y(_226_) );
INVX1 INVX1_11 ( .A(_226_), .Y(_227_) );
NAND2X1 NAND2X1_77 ( .A(_63_), .B(_37_), .Y(_228_) );
NAND3X1 NAND3X1_32 ( .A(_61_), .B(_62_), .C(_32_), .Y(_229_) );
NAND3X1 NAND3X1_33 ( .A(_227_), .B(_228_), .C(_229_), .Y(_230_) );
AOI21X1 AOI21X1_15 ( .A(_61_), .B(_62_), .C(_32_), .Y(_231_) );
NOR2X1 NOR2X1_20 ( .A(_63_), .B(_37_), .Y(_232_) );
OAI21X1 OAI21X1_24 ( .A(_231_), .B(_232_), .C(_226_), .Y(_233_) );
XNOR2X1 XNOR2X1_14 ( .A(data_in[1]), .B(_539__29_bF_buf0), .Y(_234_) );
XNOR2X1 XNOR2X1_15 ( .A(_234_), .B(data_in[5]), .Y(_235_) );
INVX1 INVX1_12 ( .A(_235_), .Y(_236_) );
NAND3X1 NAND3X1_34 ( .A(_230_), .B(_233_), .C(_236_), .Y(_237_) );
NOR3X1 NOR3X1_5 ( .A(_226_), .B(_231_), .C(_232_), .Y(_238_) );
AOI21X1 AOI21X1_16 ( .A(_229_), .B(_228_), .C(_227_), .Y(_239_) );
OAI21X1 OAI21X1_25 ( .A(_239_), .B(_238_), .C(_235_), .Y(_240_) );
NAND3X1 NAND3X1_35 ( .A(crc_en_bF_buf4), .B(_237_), .C(_240_), .Y(_241_) );
NAND2X1 NAND2X1_78 ( .A(_225_), .B(_241_), .Y(_0__9_) );
INVX1 INVX1_13 ( .A(_539__10_), .Y(_242_) );
XOR2X1 XOR2X1_14 ( .A(data_in[0]), .B(_539__29_bF_buf3), .Y(_243_) );
OAI21X1 OAI21X1_26 ( .A(_65_), .B(_66_), .C(_243_), .Y(_244_) );
XNOR2X1 XNOR2X1_16 ( .A(data_in[0]), .B(_539__29_bF_buf2), .Y(_245_) );
OAI21X1 OAI21X1_27 ( .A(_69_), .B(_70_), .C(_245_), .Y(_246_) );
NOR2X1 NOR2X1_21 ( .A(_539__27_), .B(_59_), .Y(_247_) );
NOR2X1 NOR2X1_22 ( .A(data_in[2]), .B(_68_), .Y(_248_) );
OAI21X1 OAI21X1_28 ( .A(_247_), .B(_248_), .C(_539__2_), .Y(_249_) );
NOR2X1 NOR2X1_23 ( .A(_59_), .B(_68_), .Y(_250_) );
NOR2X1 NOR2X1_24 ( .A(data_in[2]), .B(_539__27_), .Y(_251_) );
OAI21X1 OAI21X1_29 ( .A(_251_), .B(_250_), .C(_21_), .Y(_252_) );
AOI22X1 AOI22X1_9 ( .A(_249_), .B(_252_), .C(_246_), .D(_244_), .Y(_253_) );
OAI21X1 OAI21X1_30 ( .A(_65_), .B(_66_), .C(_245_), .Y(_254_) );
OAI21X1 OAI21X1_31 ( .A(_69_), .B(_70_), .C(_243_), .Y(_255_) );
NAND2X1 NAND2X1_79 ( .A(_249_), .B(_252_), .Y(_256_) );
AOI21X1 AOI21X1_17 ( .A(_254_), .B(_255_), .C(_256_), .Y(_257_) );
OAI21X1 OAI21X1_32 ( .A(_253_), .B(_257_), .C(_189_), .Y(_258_) );
AOI22X1 AOI22X1_10 ( .A(_249_), .B(_252_), .C(_254_), .D(_255_), .Y(_259_) );
AOI21X1 AOI21X1_18 ( .A(_244_), .B(_246_), .C(_256_), .Y(_260_) );
OAI21X1 OAI21X1_33 ( .A(_259_), .B(_260_), .C(_185_), .Y(_261_) );
NAND3X1 NAND3X1_36 ( .A(crc_en_bF_buf3), .B(_258_), .C(_261_), .Y(_262_) );
OAI21X1 OAI21X1_34 ( .A(crc_en_bF_buf2), .B(_242_), .C(_262_), .Y(_0__10_) );
XNOR2X1 XNOR2X1_17 ( .A(data_in_3_bF_buf1), .B(_539__3_), .Y(_263_) );
XNOR2X1 XNOR2X1_18 ( .A(_212_), .B(_263_), .Y(_264_) );
NAND3X1 NAND3X1_37 ( .A(_208_), .B(_264_), .C(_211_), .Y(_265_) );
XOR2X1 XOR2X1_15 ( .A(_212_), .B(_263_), .Y(_266_) );
NAND3X1 NAND3X1_38 ( .A(_218_), .B(_266_), .C(_220_), .Y(_267_) );
NAND2X1 NAND2X1_80 ( .A(_265_), .B(_267_), .Y(_268_) );
NAND2X1 NAND2X1_81 ( .A(_539__11_), .B(_516__bF_buf4), .Y(_269_) );
OAI21X1 OAI21X1_35 ( .A(_516__bF_buf3), .B(_268_), .C(_269_), .Y(_0__11_) );
INVX1 INVX1_14 ( .A(_539__12_), .Y(_270_) );
XNOR2X1 XNOR2X1_19 ( .A(_539__28_bF_buf2), .B(_539__29_bF_buf1), .Y(_271_) );
OAI21X1 OAI21X1_36 ( .A(_201_), .B(_202_), .C(_271_), .Y(_272_) );
NAND2X1 NAND2X1_82 ( .A(_539__28_bF_buf1), .B(_102_), .Y(_273_) );
NAND2X1 NAND2X1_83 ( .A(_539__29_bF_buf0), .B(_60_), .Y(_274_) );
NAND2X1 NAND2X1_84 ( .A(_273_), .B(_274_), .Y(_275_) );
NAND2X1 NAND2X1_85 ( .A(_275_), .B(_206_), .Y(_276_) );
NAND2X1 NAND2X1_86 ( .A(data_in[0]), .B(data_in[1]), .Y(_277_) );
NAND2X1 NAND2X1_87 ( .A(_529_), .B(_525_), .Y(_278_) );
NAND3X1 NAND3X1_39 ( .A(data_in[6]), .B(_277_), .C(_278_), .Y(_279_) );
OAI21X1 OAI21X1_37 ( .A(_127_), .B(_126_), .C(_5_), .Y(_280_) );
NAND2X1 NAND2X1_88 ( .A(_280_), .B(_279_), .Y(_281_) );
NAND3X1 NAND3X1_40 ( .A(_272_), .B(_276_), .C(_281_), .Y(_282_) );
NAND2X1 NAND2X1_89 ( .A(_539__24_), .B(_530_), .Y(_283_) );
NAND2X1 NAND2X1_90 ( .A(_539__25_), .B(_13_), .Y(_284_) );
NAND2X1 NAND2X1_91 ( .A(_539__28_bF_buf0), .B(_539__29_bF_buf3), .Y(_285_) );
NAND2X1 NAND2X1_92 ( .A(_60_), .B(_102_), .Y(_286_) );
AOI22X1 AOI22X1_11 ( .A(_283_), .B(_284_), .C(_285_), .D(_286_), .Y(_287_) );
AOI22X1 AOI22X1_12 ( .A(_273_), .B(_274_), .C(_204_), .D(_205_), .Y(_288_) );
NOR3X1 NOR3X1_6 ( .A(data_in[6]), .B(_127_), .C(_126_), .Y(_289_) );
AOI21X1 AOI21X1_19 ( .A(_278_), .B(_277_), .C(_5_), .Y(_290_) );
OAI22X1 OAI22X1_6 ( .A(_289_), .B(_290_), .C(_287_), .D(_288_), .Y(_291_) );
NAND2X1 NAND2X1_93 ( .A(_291_), .B(_282_), .Y(_292_) );
XNOR2X1 XNOR2X1_20 ( .A(data_in[2]), .B(_539__4_), .Y(_293_) );
INVX1 INVX1_15 ( .A(_293_), .Y(_294_) );
NAND2X1 NAND2X1_94 ( .A(data_in[4]), .B(_119_), .Y(_295_) );
NAND2X1 NAND2X1_95 ( .A(data_in[5]), .B(_73_), .Y(_296_) );
NAND2X1 NAND2X1_96 ( .A(_539__30_bF_buf1), .B(_29_), .Y(_297_) );
INVX2 INVX2_8 ( .A(_539__30_bF_buf0), .Y(_298_) );
NAND2X1 NAND2X1_97 ( .A(_539__26_), .B(_298_), .Y(_299_) );
AOI22X1 AOI22X1_13 ( .A(_295_), .B(_296_), .C(_297_), .D(_299_), .Y(_300_) );
NAND2X1 NAND2X1_98 ( .A(data_in[4]), .B(data_in[5]), .Y(_301_) );
NAND2X1 NAND2X1_99 ( .A(_73_), .B(_119_), .Y(_302_) );
NAND2X1 NAND2X1_100 ( .A(_539__30_bF_buf3), .B(_539__26_), .Y(_303_) );
NAND2X1 NAND2X1_101 ( .A(_298_), .B(_29_), .Y(_304_) );
AOI22X1 AOI22X1_14 ( .A(_302_), .B(_301_), .C(_303_), .D(_304_), .Y(_305_) );
OAI21X1 OAI21X1_38 ( .A(_300_), .B(_305_), .C(_294_), .Y(_306_) );
AND2X2 AND2X2_8 ( .A(data_in[4]), .B(data_in[5]), .Y(_307_) );
NOR2X1 NOR2X1_25 ( .A(data_in[4]), .B(data_in[5]), .Y(_308_) );
NOR2X1 NOR2X1_26 ( .A(_308_), .B(_307_), .Y(_309_) );
NOR2X1 NOR2X1_27 ( .A(_539__26_), .B(_298_), .Y(_310_) );
NOR2X1 NOR2X1_28 ( .A(_539__30_bF_buf2), .B(_29_), .Y(_311_) );
OAI21X1 OAI21X1_39 ( .A(_310_), .B(_311_), .C(_309_), .Y(_312_) );
INVX1 INVX1_16 ( .A(_303_), .Y(_313_) );
NOR2X1 NOR2X1_29 ( .A(_539__30_bF_buf1), .B(_539__26_), .Y(_314_) );
OAI22X1 OAI22X1_7 ( .A(_307_), .B(_308_), .C(_314_), .D(_313_), .Y(_315_) );
NAND3X1 NAND3X1_41 ( .A(_293_), .B(_315_), .C(_312_), .Y(_316_) );
AND2X2 AND2X2_9 ( .A(_316_), .B(_306_), .Y(_317_) );
NAND2X1 NAND2X1_102 ( .A(_292_), .B(_317_), .Y(_318_) );
NAND2X1 NAND2X1_103 ( .A(_306_), .B(_316_), .Y(_319_) );
NAND3X1 NAND3X1_42 ( .A(_282_), .B(_291_), .C(_319_), .Y(_320_) );
NAND3X1 NAND3X1_43 ( .A(crc_en_bF_buf1), .B(_320_), .C(_318_), .Y(_321_) );
OAI21X1 OAI21X1_40 ( .A(crc_en_bF_buf0), .B(_270_), .C(_321_), .Y(_0__12_) );
NAND2X1 NAND2X1_104 ( .A(_539__13_), .B(_516__bF_buf2), .Y(_322_) );
NAND2X1 NAND2X1_105 ( .A(data_in[1]), .B(data_in[2]), .Y(_323_) );
NAND2X1 NAND2X1_106 ( .A(_525_), .B(_59_), .Y(_324_) );
NAND2X1 NAND2X1_107 ( .A(_323_), .B(_324_), .Y(_325_) );
NAND2X1 NAND2X1_108 ( .A(_539__30_bF_buf0), .B(_530_), .Y(_326_) );
NAND2X1 NAND2X1_109 ( .A(_539__25_), .B(_298_), .Y(_327_) );
NAND2X1 NAND2X1_110 ( .A(_326_), .B(_327_), .Y(_328_) );
NAND2X1 NAND2X1_111 ( .A(_325_), .B(_328_), .Y(_329_) );
NAND2X1 NAND2X1_112 ( .A(_539__30_bF_buf3), .B(_539__25_), .Y(_330_) );
NAND2X1 NAND2X1_113 ( .A(_298_), .B(_530_), .Y(_331_) );
NAND2X1 NAND2X1_114 ( .A(_330_), .B(_331_), .Y(_332_) );
NAND3X1 NAND3X1_44 ( .A(_323_), .B(_324_), .C(_332_), .Y(_333_) );
XOR2X1 XOR2X1_16 ( .A(_539__26_), .B(_539__29_bF_buf2), .Y(_334_) );
NAND3X1 NAND3X1_45 ( .A(_334_), .B(_329_), .C(_333_), .Y(_335_) );
AOI22X1 AOI22X1_15 ( .A(_326_), .B(_327_), .C(_323_), .D(_324_), .Y(_336_) );
NAND2X1 NAND2X1_115 ( .A(data_in[1]), .B(_59_), .Y(_337_) );
NAND2X1 NAND2X1_116 ( .A(data_in[2]), .B(_525_), .Y(_338_) );
AOI22X1 AOI22X1_16 ( .A(_337_), .B(_338_), .C(_330_), .D(_331_), .Y(_339_) );
INVX1 INVX1_17 ( .A(_334_), .Y(_340_) );
OAI21X1 OAI21X1_41 ( .A(_336_), .B(_339_), .C(_340_), .Y(_341_) );
NAND2X1 NAND2X1_117 ( .A(_341_), .B(_335_), .Y(_342_) );
INVX1 INVX1_18 ( .A(_539__5_), .Y(_343_) );
NAND2X1 NAND2X1_118 ( .A(_539__31_bF_buf3), .B(data_in_3_bF_buf0), .Y(_344_) );
OR2X2 OR2X2_5 ( .A(_539__31_bF_buf2), .B(data_in_3_bF_buf3), .Y(_345_) );
NAND3X1 NAND3X1_46 ( .A(_343_), .B(_344_), .C(_345_), .Y(_346_) );
AND2X2 AND2X2_10 ( .A(_539__31_bF_buf1), .B(data_in_3_bF_buf2), .Y(_347_) );
NOR2X1 NOR2X1_30 ( .A(_539__31_bF_buf0), .B(data_in_3_bF_buf1), .Y(_348_) );
OAI21X1 OAI21X1_42 ( .A(_348_), .B(_347_), .C(_539__5_), .Y(_349_) );
NAND2X1 NAND2X1_119 ( .A(_349_), .B(_346_), .Y(_350_) );
NOR2X1 NOR2X1_31 ( .A(_125_), .B(_124_), .Y(_351_) );
NAND2X1 NAND2X1_120 ( .A(data_in[7]), .B(_68_), .Y(_352_) );
NAND2X1 NAND2X1_121 ( .A(_539__27_), .B(_6_), .Y(_353_) );
NAND3X1 NAND3X1_47 ( .A(_352_), .B(_353_), .C(_351_), .Y(_354_) );
XOR2X1 XOR2X1_17 ( .A(data_in[7]), .B(_539__27_), .Y(_355_) );
OAI21X1 OAI21X1_43 ( .A(_124_), .B(_125_), .C(_355_), .Y(_356_) );
NAND3X1 NAND3X1_48 ( .A(_356_), .B(_350_), .C(_354_), .Y(_357_) );
AND2X2 AND2X2_11 ( .A(_346_), .B(_349_), .Y(_358_) );
NAND2X1 NAND2X1_122 ( .A(data_in[6]), .B(_119_), .Y(_359_) );
NAND2X1 NAND2X1_123 ( .A(data_in[5]), .B(_5_), .Y(_360_) );
AOI21X1 AOI21X1_20 ( .A(_359_), .B(_360_), .C(_355_), .Y(_361_) );
AOI21X1 AOI21X1_21 ( .A(_352_), .B(_353_), .C(_351_), .Y(_362_) );
OAI21X1 OAI21X1_44 ( .A(_362_), .B(_361_), .C(_358_), .Y(_363_) );
NAND2X1 NAND2X1_124 ( .A(_357_), .B(_363_), .Y(_364_) );
NOR2X1 NOR2X1_32 ( .A(_342_), .B(_364_), .Y(_365_) );
AND2X2 AND2X2_12 ( .A(_335_), .B(_341_), .Y(_366_) );
AND2X2 AND2X2_13 ( .A(_363_), .B(_357_), .Y(_367_) );
OAI21X1 OAI21X1_45 ( .A(_366_), .B(_367_), .C(crc_en_bF_buf4), .Y(_368_) );
OAI21X1 OAI21X1_46 ( .A(_365_), .B(_368_), .C(_322_), .Y(_0__13_) );
NAND2X1 NAND2X1_125 ( .A(_539__14_), .B(_516__bF_buf1), .Y(_369_) );
XOR2X1 XOR2X1_18 ( .A(_539__31_bF_buf3), .B(_539__26_), .Y(_370_) );
OAI21X1 OAI21X1_47 ( .A(_247_), .B(_248_), .C(_18_), .Y(_371_) );
OAI21X1 OAI21X1_48 ( .A(_250_), .B(_251_), .C(_8_), .Y(_372_) );
NAND3X1 NAND3X1_49 ( .A(_370_), .B(_371_), .C(_372_), .Y(_373_) );
INVX1 INVX1_19 ( .A(_373_), .Y(_374_) );
AOI21X1 AOI21X1_22 ( .A(_372_), .B(_371_), .C(_370_), .Y(_375_) );
NOR2X1 NOR2X1_33 ( .A(_133_), .B(_132_), .Y(_376_) );
XOR2X1 XOR2X1_19 ( .A(_539__28_bF_buf3), .B(_539__6_), .Y(_377_) );
NAND2X1 NAND2X1_126 ( .A(_539__30_bF_buf2), .B(_377_), .Y(_378_) );
NOR2X1 NOR2X1_34 ( .A(_539__28_bF_buf2), .B(_539__6_), .Y(_379_) );
INVX1 INVX1_20 ( .A(_539__6_), .Y(_380_) );
NOR2X1 NOR2X1_35 ( .A(_60_), .B(_380_), .Y(_381_) );
OAI21X1 OAI21X1_49 ( .A(_379_), .B(_381_), .C(_298_), .Y(_382_) );
AOI21X1 AOI21X1_23 ( .A(_378_), .B(_382_), .C(_376_), .Y(_383_) );
INVX1 INVX1_21 ( .A(_376_), .Y(_384_) );
NOR2X1 NOR2X1_36 ( .A(_298_), .B(_60_), .Y(_385_) );
NOR2X1 NOR2X1_37 ( .A(_539__30_bF_buf1), .B(_539__28_bF_buf1), .Y(_386_) );
OAI21X1 OAI21X1_50 ( .A(_386_), .B(_385_), .C(_539__6_), .Y(_387_) );
XOR2X1 XOR2X1_20 ( .A(_539__30_bF_buf0), .B(_539__28_bF_buf0), .Y(_388_) );
NAND2X1 NAND2X1_127 ( .A(_380_), .B(_388_), .Y(_389_) );
AOI21X1 AOI21X1_24 ( .A(_389_), .B(_387_), .C(_384_), .Y(_390_) );
OAI22X1 OAI22X1_8 ( .A(_383_), .B(_390_), .C(_375_), .D(_374_), .Y(_391_) );
INVX1 INVX1_22 ( .A(_370_), .Y(_392_) );
NAND2X1 NAND2X1_128 ( .A(_371_), .B(_372_), .Y(_393_) );
NAND2X1 NAND2X1_129 ( .A(_392_), .B(_393_), .Y(_394_) );
NAND3X1 NAND3X1_50 ( .A(_384_), .B(_382_), .C(_378_), .Y(_395_) );
NAND3X1 NAND3X1_51 ( .A(_376_), .B(_387_), .C(_389_), .Y(_396_) );
NAND2X1 NAND2X1_130 ( .A(_395_), .B(_396_), .Y(_397_) );
NAND3X1 NAND3X1_52 ( .A(_373_), .B(_394_), .C(_397_), .Y(_398_) );
NAND3X1 NAND3X1_53 ( .A(crc_en_bF_buf3), .B(_398_), .C(_391_), .Y(_399_) );
NAND2X1 NAND2X1_131 ( .A(_369_), .B(_399_), .Y(_0__14_) );
INVX1 INVX1_23 ( .A(_539__15_), .Y(_400_) );
NAND2X1 NAND2X1_132 ( .A(_100_), .B(_101_), .Y(_401_) );
XNOR2X1 XNOR2X1_21 ( .A(_539__29_bF_buf1), .B(_539__7_), .Y(_402_) );
XNOR2X1 XNOR2X1_22 ( .A(_401_), .B(_402_), .Y(_403_) );
NAND2X1 NAND2X1_133 ( .A(_344_), .B(_345_), .Y(_404_) );
NOR2X1 NOR2X1_38 ( .A(_309_), .B(_404_), .Y(_405_) );
NOR2X1 NOR2X1_39 ( .A(_348_), .B(_347_), .Y(_406_) );
AOI21X1 AOI21X1_25 ( .A(_295_), .B(_296_), .C(_406_), .Y(_407_) );
OAI21X1 OAI21X1_51 ( .A(_407_), .B(_405_), .C(data_in[7]), .Y(_408_) );
OAI21X1 OAI21X1_52 ( .A(_307_), .B(_308_), .C(_406_), .Y(_409_) );
OAI21X1 OAI21X1_53 ( .A(_347_), .B(_348_), .C(_309_), .Y(_410_) );
NAND3X1 NAND3X1_54 ( .A(_6_), .B(_410_), .C(_409_), .Y(_411_) );
NAND3X1 NAND3X1_55 ( .A(_411_), .B(_408_), .C(_403_), .Y(_412_) );
XOR2X1 XOR2X1_21 ( .A(_401_), .B(_402_), .Y(_413_) );
AOI21X1 AOI21X1_26 ( .A(_409_), .B(_410_), .C(_6_), .Y(_414_) );
INVX1 INVX1_24 ( .A(_411_), .Y(_415_) );
OAI21X1 OAI21X1_54 ( .A(_414_), .B(_415_), .C(_413_), .Y(_416_) );
NAND3X1 NAND3X1_56 ( .A(crc_en_bF_buf2), .B(_412_), .C(_416_), .Y(_417_) );
OAI21X1 OAI21X1_55 ( .A(crc_en_bF_buf1), .B(_400_), .C(_417_), .Y(_0__15_) );
XNOR2X1 XNOR2X1_23 ( .A(_539__24_), .B(_539__28_bF_buf3), .Y(_418_) );
XNOR2X1 XNOR2X1_24 ( .A(_418_), .B(_309_), .Y(_419_) );
XNOR2X1 XNOR2X1_25 ( .A(_245_), .B(_539__8_), .Y(_420_) );
XNOR2X1 XNOR2X1_26 ( .A(_419_), .B(_420_), .Y(_421_) );
NAND2X1 NAND2X1_134 ( .A(_539__16_), .B(_516__bF_buf0), .Y(_422_) );
OAI21X1 OAI21X1_56 ( .A(_516__bF_buf5), .B(_421_), .C(_422_), .Y(_0__16_) );
XNOR2X1 XNOR2X1_27 ( .A(_234_), .B(_539__9_), .Y(_423_) );
XNOR2X1 XNOR2X1_28 ( .A(_332_), .B(_351_), .Y(_424_) );
XNOR2X1 XNOR2X1_29 ( .A(_424_), .B(_423_), .Y(_425_) );
NAND2X1 NAND2X1_135 ( .A(_539__17_), .B(_516__bF_buf4), .Y(_426_) );
OAI21X1 OAI21X1_57 ( .A(_516__bF_buf3), .B(_425_), .C(_426_), .Y(_0__17_) );
XNOR2X1 XNOR2X1_30 ( .A(_22_), .B(_539__10_), .Y(_427_) );
XNOR2X1 XNOR2X1_31 ( .A(data_in[7]), .B(_539__31_bF_buf2), .Y(_428_) );
XOR2X1 XOR2X1_22 ( .A(_428_), .B(_517_), .Y(_429_) );
XNOR2X1 XNOR2X1_32 ( .A(_429_), .B(_427_), .Y(_430_) );
NAND2X1 NAND2X1_136 ( .A(_539__18_), .B(_516__bF_buf2), .Y(_431_) );
OAI21X1 OAI21X1_58 ( .A(_516__bF_buf1), .B(_430_), .C(_431_), .Y(_0__18_) );
XNOR2X1 XNOR2X1_33 ( .A(_428_), .B(data_in_3_bF_buf0), .Y(_432_) );
XOR2X1 XOR2X1_23 ( .A(_539__27_), .B(_539__11_), .Y(_433_) );
XNOR2X1 XNOR2X1_34 ( .A(_432_), .B(_433_), .Y(_434_) );
NAND2X1 NAND2X1_137 ( .A(_539__19_), .B(_516__bF_buf0), .Y(_435_) );
OAI21X1 OAI21X1_59 ( .A(_516__bF_buf5), .B(_434_), .C(_435_), .Y(_0__19_) );
XNOR2X1 XNOR2X1_35 ( .A(_539__28_bF_buf2), .B(_539__12_), .Y(_436_) );
XNOR2X1 XNOR2X1_36 ( .A(_436_), .B(_73_), .Y(_437_) );
NAND2X1 NAND2X1_138 ( .A(_539__20_), .B(_516__bF_buf4), .Y(_438_) );
OAI21X1 OAI21X1_60 ( .A(_516__bF_buf3), .B(_437_), .C(_438_), .Y(_0__20_) );
XNOR2X1 XNOR2X1_37 ( .A(_539__29_bF_buf0), .B(_539__13_), .Y(_439_) );
XNOR2X1 XNOR2X1_38 ( .A(_439_), .B(_119_), .Y(_440_) );
NAND2X1 NAND2X1_139 ( .A(_539__21_), .B(_516__bF_buf2), .Y(_441_) );
OAI21X1 OAI21X1_61 ( .A(_516__bF_buf1), .B(_440_), .C(_441_), .Y(_0__21_) );
XOR2X1 XOR2X1_24 ( .A(_518_), .B(_539__14_), .Y(_442_) );
NAND2X1 NAND2X1_140 ( .A(_539__22_), .B(_516__bF_buf0), .Y(_443_) );
OAI21X1 OAI21X1_62 ( .A(_516__bF_buf5), .B(_442_), .C(_443_), .Y(_0__22_) );
INVX1 INVX1_25 ( .A(_539__23_), .Y(_444_) );
NAND2X1 NAND2X1_141 ( .A(_539__15_), .B(_532_), .Y(_445_) );
NAND2X1 NAND2X1_142 ( .A(_400_), .B(_535_), .Y(_446_) );
NAND3X1 NAND3X1_57 ( .A(_5_), .B(_445_), .C(_446_), .Y(_447_) );
NAND2X1 NAND2X1_143 ( .A(_539__15_), .B(_535_), .Y(_448_) );
NAND2X1 NAND2X1_144 ( .A(_400_), .B(_532_), .Y(_449_) );
NAND3X1 NAND3X1_58 ( .A(data_in[6]), .B(_449_), .C(_448_), .Y(_450_) );
NAND3X1 NAND3X1_59 ( .A(_538_), .B(_447_), .C(_450_), .Y(_451_) );
AOI21X1 AOI21X1_27 ( .A(_448_), .B(_449_), .C(data_in[6]), .Y(_452_) );
AOI21X1 AOI21X1_28 ( .A(_446_), .B(_445_), .C(_5_), .Y(_453_) );
OAI21X1 OAI21X1_63 ( .A(_452_), .B(_453_), .C(_16_), .Y(_454_) );
NAND3X1 NAND3X1_60 ( .A(crc_en_bF_buf0), .B(_451_), .C(_454_), .Y(_455_) );
OAI21X1 OAI21X1_64 ( .A(crc_en_bF_buf4), .B(_444_), .C(_455_), .Y(_0__23_) );
XNOR2X1 XNOR2X1_39 ( .A(_539__26_), .B(_539__16_), .Y(_456_) );
XNOR2X1 XNOR2X1_40 ( .A(_456_), .B(_525_), .Y(_457_) );
XNOR2X1 XNOR2X1_41 ( .A(data_in[7]), .B(data_in[2]), .Y(_458_) );
XNOR2X1 XNOR2X1_42 ( .A(_539__25_), .B(_539__31_bF_buf1), .Y(_459_) );
XNOR2X1 XNOR2X1_43 ( .A(_458_), .B(_459_), .Y(_460_) );
XNOR2X1 XNOR2X1_44 ( .A(_460_), .B(_457_), .Y(_461_) );
NAND2X1 NAND2X1_145 ( .A(_539__24_), .B(_516__bF_buf4), .Y(_462_) );
OAI21X1 OAI21X1_65 ( .A(_516__bF_buf3), .B(_461_), .C(_462_), .Y(_0__24_) );
XNOR2X1 XNOR2X1_45 ( .A(_539__27_), .B(data_in_3_bF_buf3), .Y(_463_) );
XNOR2X1 XNOR2X1_46 ( .A(_463_), .B(_539__17_), .Y(_464_) );
XOR2X1 XOR2X1_25 ( .A(_464_), .B(_22_), .Y(_465_) );
NAND2X1 NAND2X1_146 ( .A(_539__25_), .B(_516__bF_buf2), .Y(_466_) );
OAI21X1 OAI21X1_66 ( .A(_516__bF_buf1), .B(_465_), .C(_466_), .Y(_0__25_) );
NAND2X1 NAND2X1_147 ( .A(_526_), .B(_83_), .Y(_467_) );
OAI21X1 OAI21X1_67 ( .A(_522_), .B(_523_), .C(_86_), .Y(_468_) );
NAND3X1 NAND3X1_61 ( .A(_200_), .B(_468_), .C(_467_), .Y(_469_) );
AND2X2 AND2X2_14 ( .A(_83_), .B(_526_), .Y(_470_) );
NOR2X1 NOR2X1_40 ( .A(_526_), .B(_83_), .Y(_471_) );
OAI21X1 OAI21X1_68 ( .A(_471_), .B(_470_), .C(_209_), .Y(_472_) );
XNOR2X1 XNOR2X1_47 ( .A(_463_), .B(_539__18_), .Y(_473_) );
INVX1 INVX1_26 ( .A(_473_), .Y(_474_) );
NAND3X1 NAND3X1_62 ( .A(_469_), .B(_474_), .C(_472_), .Y(_475_) );
NAND2X1 NAND2X1_148 ( .A(_526_), .B(_200_), .Y(_476_) );
OAI21X1 OAI21X1_69 ( .A(_522_), .B(_523_), .C(_209_), .Y(_477_) );
NAND3X1 NAND3X1_63 ( .A(_86_), .B(_476_), .C(_477_), .Y(_478_) );
NAND2X1 NAND2X1_149 ( .A(_476_), .B(_477_), .Y(_479_) );
NAND2X1 NAND2X1_150 ( .A(_83_), .B(_479_), .Y(_480_) );
NAND3X1 NAND3X1_64 ( .A(_478_), .B(_473_), .C(_480_), .Y(_481_) );
NAND3X1 NAND3X1_65 ( .A(crc_en_bF_buf3), .B(_481_), .C(_475_), .Y(_482_) );
OAI21X1 OAI21X1_70 ( .A(crc_en_bF_buf2), .B(_29_), .C(_482_), .Y(_0__26_) );
NAND2X1 NAND2X1_151 ( .A(_539__19_), .B(_149_), .Y(_483_) );
INVX1 INVX1_27 ( .A(_539__19_), .Y(_484_) );
NAND2X1 NAND2X1_152 ( .A(_484_), .B(_147_), .Y(_485_) );
XNOR2X1 XNOR2X1_48 ( .A(data_in[7]), .B(data_in[5]), .Y(_486_) );
NAND3X1 NAND3X1_66 ( .A(_486_), .B(_485_), .C(_483_), .Y(_487_) );
NAND2X1 NAND2X1_153 ( .A(_539__19_), .B(_147_), .Y(_488_) );
NAND2X1 NAND2X1_154 ( .A(_484_), .B(_149_), .Y(_489_) );
INVX1 INVX1_28 ( .A(_486_), .Y(_490_) );
NAND3X1 NAND3X1_67 ( .A(_490_), .B(_488_), .C(_489_), .Y(_491_) );
XNOR2X1 XNOR2X1_49 ( .A(_539__25_), .B(data_in[1]), .Y(_492_) );
XOR2X1 XOR2X1_26 ( .A(_539__28_bF_buf1), .B(data_in[4]), .Y(_493_) );
XNOR2X1 XNOR2X1_50 ( .A(_493_), .B(_492_), .Y(_494_) );
AOI21X1 AOI21X1_29 ( .A(_487_), .B(_491_), .C(_494_), .Y(_495_) );
NAND3X1 NAND3X1_68 ( .A(_486_), .B(_488_), .C(_489_), .Y(_496_) );
NAND3X1 NAND3X1_69 ( .A(_490_), .B(_485_), .C(_483_), .Y(_497_) );
XOR2X1 XOR2X1_27 ( .A(_493_), .B(_492_), .Y(_498_) );
AOI21X1 AOI21X1_30 ( .A(_496_), .B(_497_), .C(_498_), .Y(_499_) );
OAI21X1 OAI21X1_71 ( .A(_495_), .B(_499_), .C(crc_en_bF_buf1), .Y(_500_) );
OAI21X1 OAI21X1_72 ( .A(crc_en_bF_buf0), .B(_68_), .C(_500_), .Y(_0__27_) );
XNOR2X1 XNOR2X1_51 ( .A(_182_), .B(_539__20_), .Y(_501_) );
NAND2X1 NAND2X1_155 ( .A(_297_), .B(_299_), .Y(_502_) );
XNOR2X1 XNOR2X1_52 ( .A(_502_), .B(_351_), .Y(_503_) );
OR2X2 OR2X2_6 ( .A(_503_), .B(_501_), .Y(_504_) );
NAND2X1 NAND2X1_156 ( .A(_501_), .B(_503_), .Y(_505_) );
NAND3X1 NAND3X1_70 ( .A(crc_en_bF_buf4), .B(_505_), .C(_504_), .Y(_506_) );
OAI21X1 OAI21X1_73 ( .A(crc_en_bF_buf3), .B(_60_), .C(_506_), .Y(_0__28_) );
XNOR2X1 XNOR2X1_53 ( .A(_463_), .B(_539__21_), .Y(_507_) );
XNOR2X1 XNOR2X1_54 ( .A(_429_), .B(_507_), .Y(_508_) );
NAND2X1 NAND2X1_157 ( .A(_539__29_bF_buf3), .B(_516__bF_buf0), .Y(_509_) );
OAI21X1 OAI21X1_74 ( .A(_516__bF_buf5), .B(_508_), .C(_509_), .Y(_0__29_) );
XNOR2X1 XNOR2X1_55 ( .A(_493_), .B(_539__22_), .Y(_510_) );
XNOR2X1 XNOR2X1_56 ( .A(_510_), .B(_428_), .Y(_511_) );
NAND2X1 NAND2X1_158 ( .A(_539__30_bF_buf3), .B(_516__bF_buf4), .Y(_512_) );
OAI21X1 OAI21X1_75 ( .A(_516__bF_buf3), .B(_511_), .C(_512_), .Y(_0__30_) );
XNOR2X1 XNOR2X1_57 ( .A(_539__29_bF_buf2), .B(_539__23_), .Y(_513_) );
XNOR2X1 XNOR2X1_58 ( .A(_513_), .B(_119_), .Y(_514_) );
NAND2X1 NAND2X1_159 ( .A(_539__31_bF_buf0), .B(_516__bF_buf2), .Y(_515_) );
OAI21X1 OAI21X1_76 ( .A(_516__bF_buf1), .B(_514_), .C(_515_), .Y(_0__31_) );
INVX8 INVX8_1 ( .A(rst), .Y(_540_) );
INVX8 INVX8_2 ( .A(crc_en_bF_buf2), .Y(_516_) );
XNOR2X1 XNOR2X1_59 ( .A(data_in[6]), .B(_539__30_bF_buf2), .Y(_517_) );
XNOR2X1 XNOR2X1_60 ( .A(_539__24_), .B(data_in[0]), .Y(_518_) );
XNOR2X1 XNOR2X1_61 ( .A(_517_), .B(_518_), .Y(_519_) );
NAND2X1 NAND2X1_160 ( .A(_539__0_), .B(_516__bF_buf0), .Y(_520_) );
OAI21X1 OAI21X1_77 ( .A(_516__bF_buf5), .B(_519_), .C(_520_), .Y(_0__0_) );
INVX1 INVX1_29 ( .A(_539__1_), .Y(_521_) );
NOR2X1 NOR2X1_41 ( .A(_539__30_bF_buf1), .B(_539__24_), .Y(_522_) );
AND2X2 AND2X2_15 ( .A(_539__30_bF_buf0), .B(_539__24_), .Y(_523_) );
OAI21X1 OAI21X1_78 ( .A(_522_), .B(_523_), .C(data_in[1]), .Y(_524_) );
INVX2 INVX2_9 ( .A(data_in[1]), .Y(_525_) );
NOR2X1 NOR2X1_42 ( .A(_522_), .B(_523_), .Y(_526_) );
NAND2X1 NAND2X1_161 ( .A(_525_), .B(_526_), .Y(_527_) );
NAND2X1 NAND2X1_162 ( .A(data_in[0]), .B(_539__25_), .Y(_528_) );
INVX1 INVX1_30 ( .A(data_in[0]), .Y(_529_) );
INVX4 INVX4_3 ( .A(_539__25_), .Y(_530_) );
NAND2X1 NAND2X1_163 ( .A(_529_), .B(_530_), .Y(_531_) );
NAND2X1 NAND2X1_164 ( .A(_528_), .B(_531_), .Y(_532_) );
NAND2X1 NAND2X1_165 ( .A(_539__31_bF_buf3), .B(_532_), .Y(_533_) );
INVX1 INVX1_31 ( .A(_539__31_bF_buf2), .Y(_534_) );
AND2X2 AND2X2_16 ( .A(_531_), .B(_528_), .Y(_535_) );
NAND2X1 NAND2X1_166 ( .A(_534_), .B(_535_), .Y(_536_) );
endmodule
