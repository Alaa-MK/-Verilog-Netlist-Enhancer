module sha1_core ( gnd, vdd, clk, reset_n, init, next, block, ready, digest, digest_valid);

input gnd, vdd;
input clk;
input reset_n;
input init;
input next;
output ready;
output digest_valid;
input [511:0] block;
output [159:0] digest;

BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf8) );
BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf7) );
BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf6) );
BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf5) );
BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf4) );
BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf3) );
BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf2) );
BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf1) );
BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_hier0_bF_buf0) );
BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf7) );
BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf6) );
BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf5) );
BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf4) );
BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf3) );
BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf2) );
BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf1) );
BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(_4548_), .Y(_4548__hier0_bF_buf0) );
BUFX4 BUFX4_18 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf7) );
BUFX4 BUFX4_19 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf6) );
BUFX4 BUFX4_20 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf5) );
BUFX4 BUFX4_21 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf4) );
BUFX4 BUFX4_22 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf3) );
BUFX4 BUFX4_23 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf2) );
BUFX4 BUFX4_24 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf1) );
BUFX4 BUFX4_25 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst), .Y(round_ctr_rst_hier0_bF_buf0) );
BUFX4 BUFX4_26 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf7) );
BUFX4 BUFX4_27 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf6) );
BUFX4 BUFX4_28 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf5) );
BUFX4 BUFX4_29 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf4) );
BUFX4 BUFX4_30 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf3) );
BUFX4 BUFX4_31 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf2) );
BUFX4 BUFX4_32 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf1) );
BUFX4 BUFX4_33 ( .gnd(gnd), .vdd(vdd), .A(_4547_), .Y(_4547__hier0_bF_buf0) );
BUFX4 BUFX4_34 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf8) );
BUFX4 BUFX4_35 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf7) );
BUFX4 BUFX4_36 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf6) );
BUFX4 BUFX4_37 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf5) );
BUFX4 BUFX4_38 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf4) );
BUFX4 BUFX4_39 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf3) );
BUFX4 BUFX4_40 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf2) );
BUFX4 BUFX4_41 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf1) );
BUFX4 BUFX4_42 ( .gnd(gnd), .vdd(vdd), .A(reset_n), .Y(reset_n_hier0_bF_buf0) );
BUFX4 BUFX4_43 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf11) );
BUFX4 BUFX4_44 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf10) );
BUFX4 BUFX4_45 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf9) );
BUFX4 BUFX4_46 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf8) );
BUFX4 BUFX4_47 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf7) );
BUFX4 BUFX4_48 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf6) );
BUFX4 BUFX4_49 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf5) );
BUFX4 BUFX4_50 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf4) );
BUFX4 BUFX4_51 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf3) );
BUFX4 BUFX4_52 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf2) );
BUFX4 BUFX4_53 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf1) );
BUFX4 BUFX4_54 ( .gnd(gnd), .vdd(vdd), .A(_3432_), .Y(_3432__bF_buf0) );
BUFX4 BUFX4_55 ( .gnd(gnd), .vdd(vdd), .A(_3717_), .Y(_3717__bF_buf4) );
BUFX4 BUFX4_56 ( .gnd(gnd), .vdd(vdd), .A(_3717_), .Y(_3717__bF_buf3) );
BUFX4 BUFX4_57 ( .gnd(gnd), .vdd(vdd), .A(_3717_), .Y(_3717__bF_buf2) );
BUFX4 BUFX4_58 ( .gnd(gnd), .vdd(vdd), .A(_3717_), .Y(_3717__bF_buf1) );
BUFX4 BUFX4_59 ( .gnd(gnd), .vdd(vdd), .A(_3717_), .Y(_3717__bF_buf0) );
BUFX4 BUFX4_60 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf11) );
BUFX4 BUFX4_61 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf10) );
BUFX4 BUFX4_62 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf9) );
BUFX4 BUFX4_63 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf8) );
BUFX4 BUFX4_64 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf7) );
BUFX4 BUFX4_65 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf6) );
BUFX4 BUFX4_66 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf5) );
BUFX4 BUFX4_67 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf4) );
BUFX4 BUFX4_68 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf3) );
BUFX4 BUFX4_69 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf2) );
BUFX4 BUFX4_70 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf1) );
BUFX4 BUFX4_71 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf0) );
BUFX4 BUFX4_72 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf88) );
BUFX4 BUFX4_73 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf87) );
BUFX4 BUFX4_74 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf86) );
BUFX4 BUFX4_75 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf85) );
BUFX4 BUFX4_76 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf84) );
BUFX4 BUFX4_77 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf83) );
BUFX4 BUFX4_78 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf82) );
BUFX4 BUFX4_79 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf81) );
BUFX4 BUFX4_80 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf80) );
BUFX4 BUFX4_81 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf79) );
BUFX4 BUFX4_82 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf78) );
BUFX4 BUFX4_83 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf77) );
BUFX4 BUFX4_84 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf76) );
BUFX4 BUFX4_85 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf75) );
BUFX4 BUFX4_86 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf74) );
BUFX4 BUFX4_87 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf73) );
BUFX4 BUFX4_88 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf72) );
BUFX4 BUFX4_89 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf71) );
BUFX4 BUFX4_90 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf70) );
BUFX4 BUFX4_91 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf69) );
BUFX4 BUFX4_92 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf68) );
BUFX4 BUFX4_93 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf67) );
BUFX4 BUFX4_94 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf66) );
BUFX4 BUFX4_95 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf65) );
BUFX4 BUFX4_96 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf64) );
BUFX4 BUFX4_97 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf63) );
BUFX4 BUFX4_98 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf62) );
BUFX4 BUFX4_99 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf61) );
BUFX4 BUFX4_100 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf60) );
BUFX4 BUFX4_101 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf59) );
BUFX4 BUFX4_102 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf58) );
BUFX4 BUFX4_103 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf57) );
BUFX4 BUFX4_104 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf56) );
BUFX4 BUFX4_105 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf55) );
BUFX4 BUFX4_106 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf54) );
BUFX4 BUFX4_107 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf53) );
BUFX4 BUFX4_108 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf52) );
BUFX4 BUFX4_109 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf51) );
BUFX4 BUFX4_110 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf50) );
BUFX4 BUFX4_111 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf49) );
BUFX4 BUFX4_112 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf48) );
BUFX4 BUFX4_113 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf47) );
BUFX4 BUFX4_114 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf46) );
BUFX4 BUFX4_115 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf45) );
BUFX4 BUFX4_116 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf44) );
BUFX4 BUFX4_117 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf43) );
BUFX4 BUFX4_118 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf42) );
BUFX4 BUFX4_119 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf41) );
BUFX4 BUFX4_120 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf40) );
BUFX4 BUFX4_121 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf39) );
BUFX4 BUFX4_122 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf38) );
BUFX4 BUFX4_123 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf37) );
BUFX4 BUFX4_124 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf36) );
BUFX4 BUFX4_125 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf35) );
BUFX4 BUFX4_126 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf34) );
BUFX4 BUFX4_127 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf33) );
BUFX4 BUFX4_128 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf32) );
BUFX4 BUFX4_129 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf31) );
BUFX4 BUFX4_130 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf30) );
BUFX4 BUFX4_131 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf29) );
BUFX4 BUFX4_132 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf28) );
BUFX4 BUFX4_133 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf27) );
BUFX4 BUFX4_134 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf26) );
BUFX4 BUFX4_135 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf25) );
BUFX4 BUFX4_136 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf24) );
BUFX4 BUFX4_137 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf23) );
BUFX4 BUFX4_138 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf22) );
BUFX4 BUFX4_139 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf21) );
BUFX4 BUFX4_140 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf20) );
BUFX4 BUFX4_141 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf19) );
BUFX4 BUFX4_142 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf18) );
BUFX4 BUFX4_143 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf17) );
BUFX4 BUFX4_144 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf16) );
BUFX4 BUFX4_145 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf15) );
BUFX4 BUFX4_146 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf14) );
BUFX4 BUFX4_147 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf13) );
BUFX4 BUFX4_148 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf12) );
BUFX4 BUFX4_149 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf11) );
BUFX4 BUFX4_150 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf10) );
BUFX4 BUFX4_151 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf9) );
BUFX4 BUFX4_152 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf0), .Y(clk_bF_buf8) );
BUFX4 BUFX4_153 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf8), .Y(clk_bF_buf7) );
BUFX4 BUFX4_154 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf7), .Y(clk_bF_buf6) );
BUFX4 BUFX4_155 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf6), .Y(clk_bF_buf5) );
BUFX4 BUFX4_156 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf5), .Y(clk_bF_buf4) );
BUFX4 BUFX4_157 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf4), .Y(clk_bF_buf3) );
BUFX4 BUFX4_158 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf3), .Y(clk_bF_buf2) );
BUFX4 BUFX4_159 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf2), .Y(clk_bF_buf1) );
BUFX4 BUFX4_160 ( .gnd(gnd), .vdd(vdd), .A(clk_hier0_bF_buf1), .Y(clk_bF_buf0) );
BUFX4 BUFX4_161 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .Y(_3740__bF_buf3) );
BUFX4 BUFX4_162 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .Y(_3740__bF_buf2) );
BUFX4 BUFX4_163 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .Y(_3740__bF_buf1) );
BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_3740_), .Y(_3740__bF_buf0) );
BUFX4 BUFX4_164 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .Y(_3411__bF_buf4) );
BUFX4 BUFX4_165 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .Y(_3411__bF_buf3) );
BUFX4 BUFX4_166 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .Y(_3411__bF_buf2) );
BUFX4 BUFX4_167 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .Y(_3411__bF_buf1) );
BUFX4 BUFX4_168 ( .gnd(gnd), .vdd(vdd), .A(_3411_), .Y(_3411__bF_buf0) );
BUFX4 BUFX4_169 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf10) );
BUFX4 BUFX4_170 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf9) );
BUFX4 BUFX4_171 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf8) );
BUFX4 BUFX4_172 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf7) );
BUFX4 BUFX4_173 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf6) );
BUFX4 BUFX4_174 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf5) );
BUFX4 BUFX4_175 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf4) );
BUFX4 BUFX4_176 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf3) );
BUFX4 BUFX4_177 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf2) );
BUFX4 BUFX4_178 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf1) );
BUFX4 BUFX4_179 ( .gnd(gnd), .vdd(vdd), .A(_3387_), .Y(_3387__bF_buf0) );
BUFX4 BUFX4_180 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .Y(_3405__bF_buf5) );
BUFX4 BUFX4_181 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .Y(_3405__bF_buf4) );
BUFX4 BUFX4_182 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .Y(_3405__bF_buf3) );
BUFX4 BUFX4_183 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .Y(_3405__bF_buf2) );
BUFX4 BUFX4_184 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .Y(_3405__bF_buf1) );
BUFX4 BUFX4_185 ( .gnd(gnd), .vdd(vdd), .A(_3405_), .Y(_3405__bF_buf0) );
BUFX4 BUFX4_186 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf8) );
BUFX4 BUFX4_187 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf7) );
BUFX4 BUFX4_188 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf6) );
BUFX4 BUFX4_189 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf5) );
BUFX4 BUFX4_190 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf4) );
BUFX4 BUFX4_191 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf3) );
BUFX4 BUFX4_192 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf2) );
BUFX4 BUFX4_193 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf1) );
BUFX4 BUFX4_194 ( .gnd(gnd), .vdd(vdd), .A(_2006_), .Y(_2006__bF_buf0) );
BUFX4 BUFX4_195 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf63) );
BUFX4 BUFX4_196 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf62) );
BUFX4 BUFX4_197 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf61) );
BUFX4 BUFX4_198 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf60) );
BUFX4 BUFX4_199 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf59) );
BUFX4 BUFX4_200 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf58) );
BUFX4 BUFX4_201 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf57) );
BUFX4 BUFX4_202 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf56) );
BUFX4 BUFX4_203 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf55) );
BUFX4 BUFX4_204 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf54) );
BUFX4 BUFX4_205 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf53) );
BUFX4 BUFX4_206 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf52) );
BUFX4 BUFX4_207 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf51) );
BUFX4 BUFX4_208 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf50) );
BUFX4 BUFX4_209 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf49) );
BUFX4 BUFX4_210 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf48) );
BUFX4 BUFX4_211 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf47) );
BUFX4 BUFX4_212 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf46) );
BUFX4 BUFX4_213 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf45) );
BUFX4 BUFX4_214 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf44) );
BUFX4 BUFX4_215 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf43) );
BUFX4 BUFX4_216 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf42) );
BUFX4 BUFX4_217 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf41) );
BUFX4 BUFX4_218 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf40) );
BUFX4 BUFX4_219 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf39) );
BUFX4 BUFX4_220 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf38) );
BUFX4 BUFX4_221 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf37) );
BUFX4 BUFX4_222 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf36) );
BUFX4 BUFX4_223 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf35) );
BUFX4 BUFX4_224 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf34) );
BUFX4 BUFX4_225 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf33) );
BUFX4 BUFX4_226 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf32) );
BUFX4 BUFX4_227 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf31) );
BUFX4 BUFX4_228 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf30) );
BUFX4 BUFX4_229 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf29) );
BUFX4 BUFX4_230 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf28) );
BUFX4 BUFX4_231 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf27) );
BUFX4 BUFX4_232 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf26) );
BUFX4 BUFX4_233 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf25) );
BUFX4 BUFX4_234 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf24) );
BUFX4 BUFX4_235 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf23) );
BUFX4 BUFX4_236 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf22) );
BUFX4 BUFX4_237 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf21) );
BUFX4 BUFX4_238 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf20) );
BUFX4 BUFX4_239 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf19) );
BUFX4 BUFX4_240 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf18) );
BUFX4 BUFX4_241 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf17) );
BUFX4 BUFX4_242 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf16) );
BUFX4 BUFX4_243 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf15) );
BUFX4 BUFX4_244 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf14) );
BUFX4 BUFX4_245 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf13) );
BUFX4 BUFX4_246 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf12) );
BUFX4 BUFX4_247 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf11) );
BUFX4 BUFX4_248 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf10) );
BUFX4 BUFX4_249 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf9) );
BUFX4 BUFX4_250 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf8) );
BUFX4 BUFX4_251 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf7), .Y(_4548__bF_buf7) );
BUFX4 BUFX4_252 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf6), .Y(_4548__bF_buf6) );
BUFX4 BUFX4_253 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf5), .Y(_4548__bF_buf5) );
BUFX4 BUFX4_254 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf4), .Y(_4548__bF_buf4) );
BUFX4 BUFX4_255 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf3), .Y(_4548__bF_buf3) );
BUFX4 BUFX4_256 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf2), .Y(_4548__bF_buf2) );
BUFX4 BUFX4_257 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf1), .Y(_4548__bF_buf1) );
BUFX4 BUFX4_258 ( .gnd(gnd), .vdd(vdd), .A(_4548__hier0_bF_buf0), .Y(_4548__bF_buf0) );
BUFX4 BUFX4_259 ( .gnd(gnd), .vdd(vdd), .A(_3437_), .Y(_3437__bF_buf3) );
BUFX4 BUFX4_260 ( .gnd(gnd), .vdd(vdd), .A(_3437_), .Y(_3437__bF_buf2) );
BUFX4 BUFX4_261 ( .gnd(gnd), .vdd(vdd), .A(_3437_), .Y(_3437__bF_buf1) );
BUFX4 BUFX4_262 ( .gnd(gnd), .vdd(vdd), .A(_3437_), .Y(_3437__bF_buf0) );
BUFX4 BUFX4_263 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .Y(_3722__bF_buf3) );
BUFX4 BUFX4_264 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .Y(_3722__bF_buf2) );
BUFX4 BUFX4_265 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .Y(_3722__bF_buf1) );
BUFX4 BUFX4_266 ( .gnd(gnd), .vdd(vdd), .A(_3722_), .Y(_3722__bF_buf0) );
BUFX4 BUFX4_267 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf7) );
BUFX4 BUFX4_268 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf6) );
BUFX4 BUFX4_269 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf5) );
BUFX4 BUFX4_270 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf4) );
BUFX4 BUFX4_271 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf3) );
BUFX4 BUFX4_272 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf2) );
BUFX4 BUFX4_273 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf1) );
BUFX4 BUFX4_274 ( .gnd(gnd), .vdd(vdd), .A(_3431_), .Y(_3431__bF_buf0) );
BUFX4 BUFX4_275 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .Y(_3692__bF_buf4) );
BUFX4 BUFX4_276 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .Y(_3692__bF_buf3) );
BUFX4 BUFX4_277 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .Y(_3692__bF_buf2) );
BUFX4 BUFX4_278 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .Y(_3692__bF_buf1) );
BUFX4 BUFX4_279 ( .gnd(gnd), .vdd(vdd), .A(_3692_), .Y(_3692__bF_buf0) );
BUFX4 BUFX4_280 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .Y(_3748__bF_buf4) );
BUFX4 BUFX4_281 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .Y(_3748__bF_buf3) );
BUFX4 BUFX4_282 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .Y(_3748__bF_buf2) );
BUFX4 BUFX4_283 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .Y(_3748__bF_buf1) );
BUFX4 BUFX4_284 ( .gnd(gnd), .vdd(vdd), .A(_3748_), .Y(_3748__bF_buf0) );
BUFX4 BUFX4_285 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .Y(_3710__bF_buf4) );
BUFX4 BUFX4_286 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .Y(_3710__bF_buf3) );
BUFX4 BUFX4_287 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .Y(_3710__bF_buf2) );
BUFX4 BUFX4_288 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .Y(_3710__bF_buf1) );
BUFX4 BUFX4_289 ( .gnd(gnd), .vdd(vdd), .A(_3710_), .Y(_3710__bF_buf0) );
BUFX4 BUFX4_290 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .Y(_3745__bF_buf4) );
BUFX4 BUFX4_291 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .Y(_3745__bF_buf3) );
BUFX4 BUFX4_292 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .Y(_3745__bF_buf2) );
BUFX4 BUFX4_293 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .Y(_3745__bF_buf1) );
BUFX4 BUFX4_294 ( .gnd(gnd), .vdd(vdd), .A(_3745_), .Y(_3745__bF_buf0) );
BUFX4 BUFX4_295 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .Y(_3451__bF_buf4) );
BUFX4 BUFX4_296 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .Y(_3451__bF_buf3) );
BUFX4 BUFX4_297 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .Y(_3451__bF_buf2) );
BUFX4 BUFX4_298 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .Y(_3451__bF_buf1) );
BUFX4 BUFX4_299 ( .gnd(gnd), .vdd(vdd), .A(_3451_), .Y(_3451__bF_buf0) );
BUFX4 BUFX4_300 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .Y(_3736__bF_buf3) );
BUFX4 BUFX4_301 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .Y(_3736__bF_buf2) );
BUFX4 BUFX4_302 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .Y(_3736__bF_buf1) );
BUFX4 BUFX4_303 ( .gnd(gnd), .vdd(vdd), .A(_3736_), .Y(_3736__bF_buf0) );
BUFX4 BUFX4_304 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf63) );
BUFX4 BUFX4_305 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf62) );
BUFX4 BUFX4_306 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf61) );
BUFX4 BUFX4_307 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf60) );
BUFX4 BUFX4_308 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf59) );
BUFX4 BUFX4_309 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf58) );
BUFX4 BUFX4_310 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf57) );
BUFX4 BUFX4_311 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf56) );
BUFX4 BUFX4_312 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf55) );
BUFX4 BUFX4_313 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf54) );
BUFX4 BUFX4_314 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf53) );
BUFX4 BUFX4_315 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf52) );
BUFX4 BUFX4_316 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf51) );
BUFX4 BUFX4_317 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf50) );
BUFX4 BUFX4_318 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf49) );
BUFX4 BUFX4_319 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf48) );
BUFX4 BUFX4_320 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf47) );
BUFX4 BUFX4_321 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf46) );
BUFX4 BUFX4_322 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf45) );
BUFX4 BUFX4_323 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf44) );
BUFX4 BUFX4_324 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf43) );
BUFX4 BUFX4_325 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf42) );
BUFX4 BUFX4_326 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf41) );
BUFX4 BUFX4_327 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf40) );
BUFX4 BUFX4_328 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf39) );
BUFX4 BUFX4_329 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf38) );
BUFX4 BUFX4_330 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf37) );
BUFX4 BUFX4_331 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf36) );
BUFX4 BUFX4_332 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf35) );
BUFX4 BUFX4_333 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf34) );
BUFX4 BUFX4_334 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf33) );
BUFX4 BUFX4_335 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf32) );
BUFX4 BUFX4_336 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf31) );
BUFX4 BUFX4_337 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf30) );
BUFX4 BUFX4_338 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf29) );
BUFX4 BUFX4_339 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf28) );
BUFX4 BUFX4_340 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf27) );
BUFX4 BUFX4_341 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf26) );
BUFX4 BUFX4_342 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf25) );
BUFX4 BUFX4_343 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf24) );
BUFX4 BUFX4_344 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf23) );
BUFX4 BUFX4_345 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf22) );
BUFX4 BUFX4_346 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf21) );
BUFX4 BUFX4_347 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf20) );
BUFX4 BUFX4_348 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf19) );
BUFX4 BUFX4_349 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf18) );
BUFX4 BUFX4_350 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf17) );
BUFX4 BUFX4_351 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf16) );
BUFX4 BUFX4_352 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf15) );
BUFX4 BUFX4_353 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf14) );
BUFX4 BUFX4_354 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf13) );
BUFX4 BUFX4_355 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf12) );
BUFX4 BUFX4_356 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf11) );
BUFX4 BUFX4_357 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf10) );
BUFX4 BUFX4_358 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf9) );
BUFX4 BUFX4_359 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf8) );
BUFX4 BUFX4_360 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf7), .Y(round_ctr_rst_bF_buf7) );
BUFX4 BUFX4_361 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf6), .Y(round_ctr_rst_bF_buf6) );
BUFX4 BUFX4_362 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf5), .Y(round_ctr_rst_bF_buf5) );
BUFX4 BUFX4_363 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf4), .Y(round_ctr_rst_bF_buf4) );
BUFX4 BUFX4_364 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf3), .Y(round_ctr_rst_bF_buf3) );
BUFX4 BUFX4_365 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf2), .Y(round_ctr_rst_bF_buf2) );
BUFX4 BUFX4_366 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf1), .Y(round_ctr_rst_bF_buf1) );
BUFX4 BUFX4_367 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_hier0_bF_buf0), .Y(round_ctr_rst_bF_buf0) );
BUFX4 BUFX4_368 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf7) );
BUFX4 BUFX4_369 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf6) );
BUFX4 BUFX4_370 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf5) );
BUFX4 BUFX4_371 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf4) );
BUFX4 BUFX4_372 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf3) );
BUFX4 BUFX4_373 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf2) );
BUFX4 BUFX4_374 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf1) );
BUFX4 BUFX4_375 ( .gnd(gnd), .vdd(vdd), .A(_3386_), .Y(_3386__bF_buf0) );
BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .Y(_3730__bF_buf4) );
BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .Y(_3730__bF_buf3) );
BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .Y(_3730__bF_buf2) );
BUFX4 BUFX4_376 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .Y(_3730__bF_buf1) );
BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(_3730_), .Y(_3730__bF_buf0) );
BUFX4 BUFX4_377 ( .gnd(gnd), .vdd(vdd), .A(_3727_), .Y(_3727__bF_buf3) );
BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(_3727_), .Y(_3727__bF_buf2) );
BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_3727_), .Y(_3727__bF_buf1) );
BUFX4 BUFX4_378 ( .gnd(gnd), .vdd(vdd), .A(_3727_), .Y(_3727__bF_buf0) );
BUFX4 BUFX4_379 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf11) );
BUFX4 BUFX4_380 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf10) );
BUFX4 BUFX4_381 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf9) );
BUFX4 BUFX4_382 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf8) );
BUFX4 BUFX4_383 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf7) );
BUFX4 BUFX4_384 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf6) );
BUFX4 BUFX4_385 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf5) );
BUFX4 BUFX4_386 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf4) );
BUFX4 BUFX4_387 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf3) );
BUFX4 BUFX4_388 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf2) );
BUFX4 BUFX4_389 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf1) );
BUFX4 BUFX4_390 ( .gnd(gnd), .vdd(vdd), .A(_2005_), .Y(_2005__bF_buf0) );
BUFX4 BUFX4_391 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf63) );
BUFX4 BUFX4_392 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf62) );
BUFX4 BUFX4_393 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf61) );
BUFX4 BUFX4_394 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf60) );
BUFX4 BUFX4_395 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf59) );
BUFX4 BUFX4_396 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf58) );
BUFX4 BUFX4_397 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf57) );
BUFX4 BUFX4_398 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf56) );
BUFX4 BUFX4_399 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf55) );
BUFX4 BUFX4_400 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf54) );
BUFX4 BUFX4_401 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf53) );
BUFX4 BUFX4_402 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf52) );
BUFX4 BUFX4_403 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf51) );
BUFX4 BUFX4_404 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf50) );
BUFX4 BUFX4_405 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf49) );
BUFX4 BUFX4_406 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf48) );
BUFX4 BUFX4_407 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf47) );
BUFX4 BUFX4_408 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf46) );
BUFX4 BUFX4_409 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf45) );
BUFX4 BUFX4_410 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf44) );
BUFX4 BUFX4_411 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf43) );
BUFX4 BUFX4_412 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf42) );
BUFX4 BUFX4_413 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf41) );
BUFX4 BUFX4_414 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf40) );
BUFX4 BUFX4_415 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf39) );
BUFX4 BUFX4_416 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf38) );
BUFX4 BUFX4_417 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf37) );
BUFX4 BUFX4_418 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf36) );
BUFX4 BUFX4_419 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf35) );
BUFX4 BUFX4_420 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf34) );
BUFX4 BUFX4_421 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf33) );
BUFX4 BUFX4_422 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf32) );
BUFX4 BUFX4_423 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf31) );
BUFX4 BUFX4_424 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf30) );
BUFX4 BUFX4_425 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf29) );
BUFX4 BUFX4_426 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf28) );
BUFX4 BUFX4_427 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf27) );
BUFX4 BUFX4_428 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf26) );
BUFX4 BUFX4_429 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf25) );
BUFX4 BUFX4_430 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf24) );
BUFX4 BUFX4_431 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf23) );
BUFX4 BUFX4_432 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf22) );
BUFX4 BUFX4_433 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf21) );
BUFX4 BUFX4_434 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf20) );
BUFX4 BUFX4_435 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf19) );
BUFX4 BUFX4_436 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf18) );
BUFX4 BUFX4_437 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf17) );
BUFX4 BUFX4_438 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf16) );
BUFX4 BUFX4_439 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf15) );
BUFX4 BUFX4_440 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf14) );
BUFX4 BUFX4_441 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf13) );
BUFX4 BUFX4_442 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf12) );
BUFX4 BUFX4_443 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf11) );
BUFX4 BUFX4_444 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf10) );
BUFX4 BUFX4_445 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf9) );
BUFX4 BUFX4_446 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf8) );
BUFX4 BUFX4_447 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf7), .Y(_4547__bF_buf7) );
BUFX4 BUFX4_448 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf6), .Y(_4547__bF_buf6) );
BUFX4 BUFX4_449 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf5), .Y(_4547__bF_buf5) );
BUFX4 BUFX4_450 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf4), .Y(_4547__bF_buf4) );
BUFX4 BUFX4_451 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf3), .Y(_4547__bF_buf3) );
BUFX4 BUFX4_452 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf2), .Y(_4547__bF_buf2) );
BUFX4 BUFX4_453 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf1), .Y(_4547__bF_buf1) );
BUFX4 BUFX4_454 ( .gnd(gnd), .vdd(vdd), .A(_4547__hier0_bF_buf0), .Y(_4547__bF_buf0) );
BUFX4 BUFX4_455 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .Y(_3474__bF_buf4) );
BUFX4 BUFX4_456 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .Y(_3474__bF_buf3) );
BUFX4 BUFX4_457 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .Y(_3474__bF_buf2) );
BUFX4 BUFX4_458 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .Y(_3474__bF_buf1) );
BUFX4 BUFX4_459 ( .gnd(gnd), .vdd(vdd), .A(_3474_), .Y(_3474__bF_buf0) );
BUFX4 BUFX4_460 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf88) );
BUFX4 BUFX4_461 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf87) );
BUFX4 BUFX4_462 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf86) );
BUFX4 BUFX4_463 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf85) );
BUFX4 BUFX4_464 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf84) );
BUFX4 BUFX4_465 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf83) );
BUFX4 BUFX4_466 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf82) );
BUFX4 BUFX4_467 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf81) );
BUFX4 BUFX4_468 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf80) );
BUFX4 BUFX4_469 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf79) );
BUFX4 BUFX4_470 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf78) );
BUFX4 BUFX4_471 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf77) );
BUFX4 BUFX4_472 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf76) );
BUFX4 BUFX4_473 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf75) );
BUFX4 BUFX4_474 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf74) );
BUFX4 BUFX4_475 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf73) );
BUFX4 BUFX4_476 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf72) );
BUFX4 BUFX4_477 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf71) );
BUFX4 BUFX4_478 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf70) );
BUFX4 BUFX4_479 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf69) );
BUFX4 BUFX4_480 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf68) );
BUFX4 BUFX4_481 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf67) );
BUFX4 BUFX4_482 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf66) );
BUFX4 BUFX4_483 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf65) );
BUFX4 BUFX4_484 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf64) );
BUFX4 BUFX4_485 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf63) );
BUFX4 BUFX4_486 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf62) );
BUFX4 BUFX4_487 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf61) );
BUFX4 BUFX4_488 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf60) );
BUFX4 BUFX4_489 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf59) );
BUFX4 BUFX4_490 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf58) );
BUFX4 BUFX4_491 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf57) );
BUFX4 BUFX4_492 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf56) );
BUFX4 BUFX4_493 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf55) );
BUFX4 BUFX4_494 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf54) );
BUFX4 BUFX4_495 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf53) );
BUFX4 BUFX4_496 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf52) );
BUFX4 BUFX4_497 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf51) );
BUFX4 BUFX4_498 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf50) );
BUFX4 BUFX4_499 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf49) );
BUFX4 BUFX4_500 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf48) );
BUFX4 BUFX4_501 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf47) );
BUFX4 BUFX4_502 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf46) );
BUFX4 BUFX4_503 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf45) );
BUFX4 BUFX4_504 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf44) );
BUFX4 BUFX4_505 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf43) );
BUFX4 BUFX4_506 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf42) );
BUFX4 BUFX4_507 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf41) );
BUFX4 BUFX4_508 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf40) );
BUFX4 BUFX4_509 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf39) );
BUFX4 BUFX4_510 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf38) );
BUFX4 BUFX4_511 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf37) );
BUFX4 BUFX4_512 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf36) );
BUFX4 BUFX4_513 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf35) );
BUFX4 BUFX4_514 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf34) );
BUFX4 BUFX4_515 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf33) );
BUFX4 BUFX4_516 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf32) );
BUFX4 BUFX4_517 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf31) );
BUFX4 BUFX4_518 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf30) );
BUFX4 BUFX4_519 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf29) );
BUFX4 BUFX4_520 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf28) );
BUFX4 BUFX4_521 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf27) );
BUFX4 BUFX4_522 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf26) );
BUFX4 BUFX4_523 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf25) );
BUFX4 BUFX4_524 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf24) );
BUFX4 BUFX4_525 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf23) );
BUFX4 BUFX4_526 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf22) );
BUFX4 BUFX4_527 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf21) );
BUFX4 BUFX4_528 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf20) );
BUFX4 BUFX4_529 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf19) );
BUFX4 BUFX4_530 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf18) );
BUFX4 BUFX4_531 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf17) );
BUFX4 BUFX4_532 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf16) );
BUFX4 BUFX4_533 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf15) );
BUFX4 BUFX4_534 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf14) );
BUFX4 BUFX4_535 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf13) );
BUFX4 BUFX4_536 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf12) );
BUFX4 BUFX4_537 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf11) );
BUFX4 BUFX4_538 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf10) );
BUFX4 BUFX4_539 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf9) );
BUFX4 BUFX4_540 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf8) );
BUFX4 BUFX4_541 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf7) );
BUFX4 BUFX4_542 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf6) );
BUFX4 BUFX4_543 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf5) );
BUFX4 BUFX4_544 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf4) );
BUFX4 BUFX4_545 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf3) );
BUFX4 BUFX4_546 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf2) );
BUFX4 BUFX4_547 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf1) );
BUFX4 BUFX4_548 ( .gnd(gnd), .vdd(vdd), .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf0) );
BUFX4 BUFX4_549 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf11) );
BUFX4 BUFX4_550 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf10) );
BUFX4 BUFX4_551 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf9) );
BUFX4 BUFX4_552 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf8) );
BUFX4 BUFX4_553 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf7) );
BUFX4 BUFX4_554 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf6) );
BUFX4 BUFX4_555 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf5) );
BUFX4 BUFX4_556 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf4) );
BUFX4 BUFX4_557 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf3) );
BUFX4 BUFX4_558 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf2) );
BUFX4 BUFX4_559 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf1) );
BUFX4 BUFX4_560 ( .gnd(gnd), .vdd(vdd), .A(_3433_), .Y(_3433__bF_buf0) );
BUFX4 BUFX4_561 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .Y(_3691__bF_buf4) );
BUFX4 BUFX4_562 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .Y(_3691__bF_buf3) );
BUFX4 BUFX4_563 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .Y(_3691__bF_buf2) );
BUFX4 BUFX4_564 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .Y(_3691__bF_buf1) );
BUFX4 BUFX4_565 ( .gnd(gnd), .vdd(vdd), .A(_3691_), .Y(_3691__bF_buf0) );
BUFX4 BUFX4_566 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .Y(_3747__bF_buf4) );
BUFX4 BUFX4_567 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .Y(_3747__bF_buf3) );
BUFX4 BUFX4_568 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .Y(_3747__bF_buf2) );
BUFX4 BUFX4_569 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .Y(_3747__bF_buf1) );
BUFX4 BUFX4_570 ( .gnd(gnd), .vdd(vdd), .A(_3747_), .Y(_3747__bF_buf0) );
BUFX4 BUFX4_571 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_113__bF_buf4) );
BUFX4 BUFX4_572 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_113__bF_buf3) );
BUFX4 BUFX4_573 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_113__bF_buf2) );
BUFX4 BUFX4_574 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_113__bF_buf1) );
BUFX4 BUFX4_575 ( .gnd(gnd), .vdd(vdd), .A(_113_), .Y(_113__bF_buf0) );
BUFX4 BUFX4_576 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_40__bF_buf3) );
BUFX4 BUFX4_577 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_40__bF_buf2) );
BUFX4 BUFX4_578 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_40__bF_buf1) );
BUFX4 BUFX4_579 ( .gnd(gnd), .vdd(vdd), .A(_40_), .Y(_40__bF_buf0) );
BUFX4 BUFX4_580 ( .gnd(gnd), .vdd(vdd), .A(_3706_), .Y(_3706__bF_buf3) );
BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_3706_), .Y(_3706__bF_buf2) );
BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_3706_), .Y(_3706__bF_buf1) );
BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_3706_), .Y(_3706__bF_buf0) );
BUFX4 BUFX4_581 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .Y(_3738__bF_buf4) );
BUFX4 BUFX4_582 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .Y(_3738__bF_buf3) );
BUFX4 BUFX4_583 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .Y(_3738__bF_buf2) );
BUFX4 BUFX4_584 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .Y(_3738__bF_buf1) );
BUFX4 BUFX4_585 ( .gnd(gnd), .vdd(vdd), .A(_3738_), .Y(_3738__bF_buf0) );
BUFX4 BUFX4_586 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .Y(_3700__bF_buf3) );
BUFX4 BUFX4_587 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .Y(_3700__bF_buf2) );
BUFX4 BUFX4_588 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .Y(_3700__bF_buf1) );
BUFX4 BUFX4_589 ( .gnd(gnd), .vdd(vdd), .A(_3700_), .Y(_3700__bF_buf0) );
BUFX4 BUFX4_590 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .Y(_3735__bF_buf4) );
BUFX4 BUFX4_591 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .Y(_3735__bF_buf3) );
BUFX4 BUFX4_592 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .Y(_3735__bF_buf2) );
BUFX4 BUFX4_593 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .Y(_3735__bF_buf1) );
BUFX4 BUFX4_594 ( .gnd(gnd), .vdd(vdd), .A(_3735_), .Y(_3735__bF_buf0) );
BUFX4 BUFX4_595 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .Y(_3447__bF_buf4) );
BUFX4 BUFX4_596 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .Y(_3447__bF_buf3) );
BUFX4 BUFX4_597 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .Y(_3447__bF_buf2) );
BUFX4 BUFX4_598 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .Y(_3447__bF_buf1) );
BUFX4 BUFX4_599 ( .gnd(gnd), .vdd(vdd), .A(_3447_), .Y(_3447__bF_buf0) );
BUFX4 BUFX4_600 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .Y(_3732__bF_buf4) );
BUFX4 BUFX4_601 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .Y(_3732__bF_buf3) );
BUFX4 BUFX4_602 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .Y(_3732__bF_buf2) );
BUFX4 BUFX4_603 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .Y(_3732__bF_buf1) );
BUFX4 BUFX4_604 ( .gnd(gnd), .vdd(vdd), .A(_3732_), .Y(_3732__bF_buf0) );
BUFX4 BUFX4_605 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3406__bF_buf4) );
BUFX4 BUFX4_606 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3406__bF_buf3) );
BUFX4 BUFX4_607 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3406__bF_buf2) );
BUFX4 BUFX4_608 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3406__bF_buf1) );
BUFX4 BUFX4_609 ( .gnd(gnd), .vdd(vdd), .A(_3406_), .Y(_3406__bF_buf0) );
BUFX4 BUFX4_610 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf8) );
BUFX4 BUFX4_611 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf7) );
BUFX4 BUFX4_612 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf6) );
BUFX4 BUFX4_613 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf5) );
BUFX4 BUFX4_614 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf4) );
BUFX4 BUFX4_615 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf3) );
BUFX4 BUFX4_616 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf2) );
BUFX4 BUFX4_617 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf1) );
BUFX4 BUFX4_618 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new), .Y(digest_valid_new_bF_buf0) );
XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3805_), .B(_3806_), .Y(_3807_) );
INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__3_), .Y(_3808_) );
OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(_3783_), .C(_3691__bF_buf4), .Y(_3809_) );
INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__3_), .Y(_3810_) );
NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__3_), .B(_3747__bF_buf4), .Y(_3811_) );
OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_3810_), .B(_3717__bF_buf4), .C(_3811_), .Y(_3812_) );
INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__3_), .Y(_3813_) );
INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__3_), .Y(_3814_) );
OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3814_), .B(_3764_), .C(_3813_), .D(_3763_), .Y(_3815_) );
NOR3X1 NOR3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3812_), .B(_3809_), .C(_3815_), .Y(_3816_) );
NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__3_), .B(_3710__bF_buf4), .Y(_3817_) );
NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__3_), .B(_3706__bF_buf3), .Y(_3818_) );
NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__3_), .B(_3721_), .Y(_3819_) );
NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3817_), .B(_3819_), .C(_3818_), .Y(_3820_) );
AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__3_), .B(_3745__bF_buf4), .C(w_mem_inst_w_mem_1__3_), .D(_3732__bF_buf4), .Y(_3821_) );
NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__3_), .B(_3738__bF_buf4), .Y(_3822_) );
NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__3_), .B(_3743_), .Y(_3823_) );
NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_3822_), .B(_3823_), .C(_3821_), .Y(_3824_) );
AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__3_), .B(_3736__bF_buf3), .C(w_mem_inst_w_mem_4__3_), .D(_3740__bF_buf3), .Y(_3825_) );
AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__3_), .B(_3735__bF_buf4), .C(w_mem_inst_w_mem_2__3_), .D(_3700__bF_buf3), .Y(_3826_) );
NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3825_), .B(_3826_), .Y(_3827_) );
NOR3X1 NOR3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_3820_), .B(_3827_), .C(_3824_), .Y(_3828_) );
AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf4), .B(_3807_), .C(_3816_), .D(_3828_), .Y(w_3_) );
XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__3_), .B(w_mem_inst_w_mem_13__3_), .Y(_3829_) );
XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__3_), .B(w_mem_inst_w_mem_2__3_), .Y(_3830_) );
XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3829_), .B(_3830_), .Y(_3831_) );
INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__4_), .Y(_3832_) );
INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(_3740__bF_buf2), .Y(_3833_) );
OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3832_), .B(_3833_), .C(_3691__bF_buf3), .Y(_3834_) );
INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__4_), .Y(_3835_) );
INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__4_), .Y(_3836_) );
INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf3), .Y(_3837_) );
INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(_3736__bF_buf2), .Y(_3838_) );
OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_3838_), .C(_3836_), .D(_3837_), .Y(_3839_) );
INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__4_), .Y(_3840_) );
INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__4_), .Y(_3841_) );
OAI22X1 OAI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_3756_), .C(_3840_), .D(_3763_), .Y(_3842_) );
NOR3X1 NOR3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3839_), .B(_3834_), .C(_3842_), .Y(_3843_) );
NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__4_), .B(_3732__bF_buf3), .Y(_3844_) );
NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__4_), .B(_3730__bF_buf4), .Y(_3845_) );
NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__4_), .B(_3748__bF_buf4), .Y(_3846_) );
NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3845_), .B(_3844_), .C(_3846_), .Y(_3847_) );
AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__4_), .B(_3710__bF_buf3), .C(w_mem_inst_w_mem_2__4_), .D(_3700__bF_buf2), .Y(_3848_) );
NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__4_), .B(_3745__bF_buf3), .Y(_3849_) );
NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__4_), .B(_3721_), .Y(_3850_) );
NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3849_), .B(_3850_), .C(_3848_), .Y(_3851_) );
NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__4_), .B(_3706__bF_buf2), .Y(_3852_) );
NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__4_), .B(_3747__bF_buf3), .Y(_3853_) );
AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__4_), .B(_3738__bF_buf3), .C(w_mem_inst_w_mem_13__4_), .D(_3716_), .Y(_3854_) );
NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_3853_), .B(_3854_), .C(_3852_), .Y(_3855_) );
NOR3X1 NOR3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3847_), .B(_3855_), .C(_3851_), .Y(_3856_) );
AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf3), .B(_3831_), .C(_3843_), .D(_3856_), .Y(w_4_) );
XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__4_), .B(w_mem_inst_w_mem_13__4_), .Y(_3857_) );
XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__4_), .B(w_mem_inst_w_mem_2__4_), .Y(_3858_) );
XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3857_), .B(_3858_), .Y(_3859_) );
INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__5_), .Y(_3860_) );
OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .B(_3722__bF_buf3), .C(_3691__bF_buf2), .Y(_3861_) );
INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__5_), .Y(_3862_) );
NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__5_), .B(_3747__bF_buf2), .Y(_3863_) );
OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_3862_), .B(_3763_), .C(_3863_), .Y(_3864_) );
INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__5_), .Y(_3865_) );
NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__5_), .B(_3710__bF_buf2), .Y(_3866_) );
OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3865_), .B(_3789_), .C(_3866_), .Y(_3867_) );
NOR3X1 NOR3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_3861_), .B(_3867_), .C(_3864_), .Y(_3868_) );
NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__5_), .B(_3706__bF_buf1), .Y(_3869_) );
NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__5_), .B(_3736__bF_buf1), .Y(_3870_) );
NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__5_), .B(_3716_), .Y(_3871_) );
NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3870_), .B(_3871_), .C(_3869_), .Y(_3872_) );
NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__5_), .B(_3730__bF_buf3), .Y(_3873_) );
NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__5_), .B(_3743_), .Y(_3874_) );
AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3740__bF_buf1), .B(w_mem_inst_w_mem_4__5_), .C(w_mem_inst_w_mem_10__5_), .D(_3748__bF_buf3), .Y(_3875_) );
NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3873_), .B(_3874_), .C(_3875_), .Y(_3876_) );
AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__5_), .B(_3738__bF_buf2), .C(w_mem_inst_w_mem_14__5_), .D(_3735__bF_buf2), .Y(_3877_) );
NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__5_), .B(_3700__bF_buf1), .Y(_3878_) );
NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__5_), .B(_3745__bF_buf2), .Y(_3879_) );
NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3879_), .B(_3878_), .C(_3877_), .Y(_3880_) );
NOR3X1 NOR3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3872_), .B(_3880_), .C(_3876_), .Y(_3881_) );
AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf2), .B(_3859_), .C(_3868_), .D(_3881_), .Y(w_5_) );
XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__5_), .B(w_mem_inst_w_mem_13__5_), .Y(_3882_) );
XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__5_), .B(w_mem_inst_w_mem_2__5_), .Y(_3883_) );
XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3882_), .B(_3883_), .Y(_3884_) );
INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__6_), .Y(_3885_) );
OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .B(_3837_), .C(_3691__bF_buf1), .Y(_3886_) );
INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__6_), .Y(_3887_) );
INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__6_), .Y(_3888_) );
OAI22X1 OAI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(_3888_), .B(_3838_), .C(_3887_), .D(_3763_), .Y(_3889_) );
INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__6_), .Y(_3890_) );
INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__6_), .Y(_3891_) );
OAI22X1 OAI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_3890_), .B(_3717__bF_buf3), .C(_3891_), .D(_3756_), .Y(_3892_) );
NOR3X1 NOR3X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3886_), .B(_3892_), .C(_3889_), .Y(_3893_) );
NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__6_), .B(_3732__bF_buf2), .Y(_3894_) );
NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__6_), .B(_3730__bF_buf2), .Y(_3895_) );
NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__6_), .B(_3747__bF_buf1), .Y(_3896_) );
NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3895_), .B(_3896_), .C(_3894_), .Y(_3897_) );
AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__6_), .B(_3710__bF_buf1), .C(w_mem_inst_w_mem_2__6_), .D(_3700__bF_buf0), .Y(_3898_) );
AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__6_), .B(_3745__bF_buf1), .C(w_mem_inst_w_mem_4__6_), .D(_3740__bF_buf0), .Y(_3899_) );
NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3898_), .B(_3899_), .Y(_3900_) );
NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__6_), .B(_3706__bF_buf0), .Y(_3901_) );
NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__6_), .B(_3721_), .Y(_3902_) );
AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__6_), .B(_3738__bF_buf1), .C(w_mem_inst_w_mem_10__6_), .D(_3748__bF_buf2), .Y(_3903_) );
NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3901_), .B(_3902_), .C(_3903_), .Y(_3904_) );
NOR3X1 NOR3X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3897_), .B(_3900_), .C(_3904_), .Y(_3905_) );
AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf1), .B(_3884_), .C(_3893_), .D(_3905_), .Y(w_6_) );
XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__6_), .B(w_mem_inst_w_mem_13__6_), .Y(_3906_) );
XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__6_), .B(w_mem_inst_w_mem_2__6_), .Y(_3907_) );
XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_3906_), .B(_3907_), .Y(_3908_) );
INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__7_), .Y(_3909_) );
OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3909_), .B(_3833_), .C(_3691__bF_buf0), .Y(_3910_) );
INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__7_), .Y(_3911_) );
NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__7_), .B(_3747__bF_buf0), .Y(_3912_) );
OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(_3717__bF_buf2), .C(_3912_), .Y(_3913_) );
INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__7_), .Y(_3914_) );
NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__7_), .B(_3710__bF_buf0), .Y(_3915_) );
OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_3707_), .C(_3915_), .Y(_3916_) );
NOR3X1 NOR3X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3913_), .B(_3910_), .C(_3916_), .Y(_3917_) );
NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__7_), .B(_3738__bF_buf0), .Y(_3918_) );
NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__7_), .B(_3730__bF_buf1), .Y(_3919_) );
NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__7_), .B(_3732__bF_buf1), .Y(_3920_) );
NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_3918_), .B(_3919_), .C(_3920_), .Y(_3921_) );
AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__7_), .B(_3736__bF_buf0), .C(w_mem_inst_w_mem_8__7_), .D(_3721_), .Y(_3922_) );
NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__7_), .B(_3700__bF_buf3), .Y(_3923_) );
NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__7_), .B(_3748__bF_buf1), .Y(_3924_) );
NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3923_), .B(_3924_), .C(_3922_), .Y(_3925_) );
AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__7_), .B(_3745__bF_buf0), .C(w_mem_inst_w_mem_5__7_), .D(_3743_), .Y(_3926_) );
AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__7_), .B(_3735__bF_buf1), .C(w_mem_inst_w_mem_9__7_), .D(_3727__bF_buf3), .Y(_3927_) );
NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_3926_), .B(_3927_), .Y(_3928_) );
NOR3X1 NOR3X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3921_), .B(_3928_), .C(_3925_), .Y(_3929_) );
AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf0), .B(_3908_), .C(_3917_), .D(_3929_), .Y(w_7_) );
XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__7_), .B(w_mem_inst_w_mem_13__7_), .Y(_3930_) );
XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__7_), .B(w_mem_inst_w_mem_2__7_), .Y(_3931_) );
XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_3930_), .B(_3931_), .Y(_3932_) );
INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__8_), .Y(_3933_) );
OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_3933_), .B(_3707_), .C(_3691__bF_buf4), .Y(_3934_) );
INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__8_), .Y(_3935_) );
INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__8_), .Y(_3936_) );
OAI22X1 OAI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3936_), .B(_3722__bF_buf2), .C(_3935_), .D(_3783_), .Y(_3937_) );
INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__8_), .Y(_3938_) );
INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__8_), .Y(_3939_) );
OAI22X1 OAI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3938_), .B(_3838_), .C(_3939_), .D(_3764_), .Y(_3940_) );
NOR3X1 NOR3X1_11 ( .gnd(gnd), .vdd(vdd), .A(_3940_), .B(_3934_), .C(_3937_), .Y(_3941_) );
NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__8_), .B(_3738__bF_buf4), .Y(_3942_) );
NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__8_), .B(_3745__bF_buf4), .Y(_3943_) );
NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__8_), .B(_3740__bF_buf3), .Y(_3944_) );
NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_3942_), .B(_3943_), .C(_3944_), .Y(_3945_) );
NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__8_), .B(_3727__bF_buf2), .Y(_3946_) );
NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__8_), .B(_3700__bF_buf2), .Y(_3947_) );
AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__8_), .B(_3710__bF_buf4), .C(w_mem_inst_w_mem_1__8_), .D(_3732__bF_buf0), .Y(_3948_) );
NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3946_), .B(_3947_), .C(_3948_), .Y(_3949_) );
AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(w_mem_inst_w_mem_13__8_), .C(w_mem_inst_w_mem_14__8_), .D(_3735__bF_buf0), .Y(_3950_) );
NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__8_), .B(_3747__bF_buf4), .Y(_3951_) );
NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__8_), .B(_3743_), .Y(_3952_) );
NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_3951_), .B(_3952_), .C(_3950_), .Y(_3953_) );
NOR3X1 NOR3X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3945_), .B(_3953_), .C(_3949_), .Y(_3954_) );
AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf4), .B(_3932_), .C(_3941_), .D(_3954_), .Y(w_8_) );
XNOR2X1 XNOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__8_), .B(w_mem_inst_w_mem_13__8_), .Y(_3955_) );
XNOR2X1 XNOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__8_), .B(w_mem_inst_w_mem_2__8_), .Y(_3956_) );
XNOR2X1 XNOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_3955_), .B(_3956_), .Y(_3957_) );
INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__9_), .Y(_3958_) );
OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3958_), .B(_3764_), .C(_3691__bF_buf3), .Y(_3959_) );
INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__9_), .Y(_3960_) );
INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__9_), .Y(_3961_) );
OAI22X1 OAI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_3756_), .C(_3960_), .D(_3701_), .Y(_3962_) );
INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__9_), .Y(_3963_) );
INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__9_), .Y(_3964_) );
OAI22X1 OAI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .B(_3717__bF_buf1), .C(_3963_), .D(_3722__bF_buf1), .Y(_3965_) );
NOR3X1 NOR3X1_13 ( .gnd(gnd), .vdd(vdd), .A(_3959_), .B(_3962_), .C(_3965_), .Y(_3966_) );
NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__9_), .B(_3727__bF_buf1), .Y(_3967_) );
NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__9_), .B(_3732__bF_buf4), .Y(_3968_) );
NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__9_), .B(_3740__bF_buf2), .Y(_3969_) );
NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_3968_), .B(_3969_), .C(_3967_), .Y(_3970_) );
AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf4), .B(w_mem_inst_w_mem_14__9_), .C(w_mem_inst_w_mem_7__9_), .D(_3736__bF_buf3), .Y(_3971_) );
NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__9_), .B(_3738__bF_buf3), .Y(_3972_) );
NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__9_), .B(_3706__bF_buf3), .Y(_3973_) );
NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_3972_), .B(_3973_), .C(_3971_), .Y(_3974_) );
AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3745__bF_buf3), .B(w_mem_inst_w_mem_11__9_), .C(w_mem_inst_w_mem_0__9_), .D(_3710__bF_buf3), .Y(_3975_) );
NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__9_), .B(_3747__bF_buf3), .Y(_3976_) );
NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__9_), .B(_3748__bF_buf0), .Y(_3977_) );
NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_3976_), .B(_3977_), .C(_3975_), .Y(_3978_) );
NOR3X1 NOR3X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3970_), .B(_3974_), .C(_3978_), .Y(_3979_) );
AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf3), .B(_3957_), .C(_3966_), .D(_3979_), .Y(w_9_) );
XNOR2X1 XNOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__9_), .B(w_mem_inst_w_mem_13__9_), .Y(_3980_) );
XNOR2X1 XNOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__9_), .B(w_mem_inst_w_mem_2__9_), .Y(_3981_) );
XNOR2X1 XNOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3980_), .B(_3981_), .Y(_3982_) );
INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__10_), .Y(_3983_) );
OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_3983_), .B(_3701_), .C(_3691__bF_buf2), .Y(_3984_) );
INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__10_), .Y(_3985_) );
NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__10_), .B(_3710__bF_buf2), .Y(_3986_) );
OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3985_), .B(_3756_), .C(_3986_), .Y(_3987_) );
INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__10_), .Y(_3988_) );
INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__10_), .Y(_3989_) );
OAI22X1 OAI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .B(_3717__bF_buf0), .C(_3988_), .D(_3722__bF_buf0), .Y(_3990_) );
NOR3X1 NOR3X1_15 ( .gnd(gnd), .vdd(vdd), .A(_3987_), .B(_3984_), .C(_3990_), .Y(_3991_) );
NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__10_), .B(_3727__bF_buf0), .Y(_3992_) );
NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__10_), .B(_3730__bF_buf0), .Y(_3993_) );
NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__10_), .B(_3732__bF_buf3), .Y(_3994_) );
NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_3993_), .B(_3994_), .C(_3992_), .Y(_3995_) );
AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf3), .B(w_mem_inst_w_mem_14__10_), .C(w_mem_inst_w_mem_7__10_), .D(_3736__bF_buf2), .Y(_3996_) );
NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__10_), .B(_3738__bF_buf2), .Y(_3997_) );
NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__10_), .B(_3740__bF_buf1), .Y(_3998_) );
NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3997_), .B(_3998_), .C(_3996_), .Y(_3999_) );
NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__10_), .B(_3706__bF_buf2), .Y(_4000_) );
NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__10_), .B(_3745__bF_buf2), .Y(_4001_) );
AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf2), .B(w_mem_inst_w_mem_12__10_), .C(w_mem_inst_w_mem_10__10_), .D(_3748__bF_buf4), .Y(_4002_) );
NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_4000_), .B(_4001_), .C(_4002_), .Y(_4003_) );
NOR3X1 NOR3X1_16 ( .gnd(gnd), .vdd(vdd), .A(_3995_), .B(_3999_), .C(_4003_), .Y(_4004_) );
AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf2), .B(_3982_), .C(_3991_), .D(_4004_), .Y(w_10_) );
XNOR2X1 XNOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__10_), .B(w_mem_inst_w_mem_13__10_), .Y(_4005_) );
XNOR2X1 XNOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__10_), .B(w_mem_inst_w_mem_2__10_), .Y(_4006_) );
XNOR2X1 XNOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_4005_), .B(_4006_), .Y(_4007_) );
INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__11_), .Y(_4008_) );
OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .B(_3833_), .C(_3691__bF_buf1), .Y(_4009_) );
INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__11_), .Y(_4010_) );
NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__11_), .B(_3710__bF_buf1), .Y(_4011_) );
OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_3707_), .C(_4011_), .Y(_4012_) );
INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__11_), .Y(_4013_) );
INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__11_), .Y(_4014_) );
OAI22X1 OAI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_3717__bF_buf4), .C(_4013_), .D(_3722__bF_buf3), .Y(_4015_) );
NOR3X1 NOR3X1_17 ( .gnd(gnd), .vdd(vdd), .A(_4009_), .B(_4015_), .C(_4012_), .Y(_4016_) );
NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__11_), .B(_3727__bF_buf3), .Y(_4017_) );
NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__11_), .B(_3730__bF_buf4), .Y(_4018_) );
NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__11_), .B(_3732__bF_buf2), .Y(_4019_) );
NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_4018_), .B(_4019_), .C(_4017_), .Y(_4020_) );
AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf2), .B(w_mem_inst_w_mem_14__11_), .C(w_mem_inst_w_mem_7__11_), .D(_3736__bF_buf1), .Y(_4021_) );
NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__11_), .B(_3738__bF_buf1), .Y(_4022_) );
NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__11_), .B(_3700__bF_buf1), .Y(_4023_) );
NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_4022_), .B(_4023_), .C(_4021_), .Y(_4024_) );
NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__11_), .B(_3743_), .Y(_4025_) );
NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__11_), .B(_3745__bF_buf1), .Y(_4026_) );
AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf1), .B(w_mem_inst_w_mem_12__11_), .C(w_mem_inst_w_mem_10__11_), .D(_3748__bF_buf3), .Y(_4027_) );
NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_4025_), .B(_4026_), .C(_4027_), .Y(_4028_) );
NOR3X1 NOR3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_4020_), .B(_4024_), .C(_4028_), .Y(_4029_) );
AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf1), .B(_4007_), .C(_4016_), .D(_4029_), .Y(w_11_) );
XNOR2X1 XNOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__11_), .B(w_mem_inst_w_mem_13__11_), .Y(_4030_) );
XNOR2X1 XNOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__11_), .B(w_mem_inst_w_mem_2__11_), .Y(_4031_) );
XNOR2X1 XNOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_4030_), .B(_4031_), .Y(_4032_) );
INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__12_), .Y(_4033_) );
OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .B(_3833_), .C(_3691__bF_buf0), .Y(_4034_) );
INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__12_), .Y(_4035_) );
INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__12_), .Y(_4036_) );
OAI22X1 OAI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .B(_3838_), .C(_4035_), .D(_3763_), .Y(_4037_) );
INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__12_), .Y(_4038_) );
INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__12_), .Y(_4039_) );
OAI22X1 OAI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .B(_3717__bF_buf3), .C(_4039_), .D(_3756_), .Y(_4040_) );
NOR3X1 NOR3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_4040_), .B(_4034_), .C(_4037_), .Y(_4041_) );
NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__12_), .B(_3732__bF_buf1), .Y(_4042_) );
NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__12_), .B(_3730__bF_buf3), .Y(_4043_) );
NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__12_), .B(_3747__bF_buf0), .Y(_4044_) );
NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_4043_), .B(_4044_), .C(_4042_), .Y(_4045_) );
NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__12_), .B(_3710__bF_buf0), .Y(_4046_) );
NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__12_), .B(_3700__bF_buf0), .Y(_4047_) );
AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf1), .B(w_mem_inst_w_mem_14__12_), .C(w_mem_inst_w_mem_11__12_), .D(_3745__bF_buf0), .Y(_4048_) );
NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_4046_), .B(_4047_), .C(_4048_), .Y(_4049_) );
NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__12_), .B(_3706__bF_buf1), .Y(_4050_) );
NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__12_), .B(_3721_), .Y(_4051_) );
AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__12_), .B(_3738__bF_buf0), .C(w_mem_inst_w_mem_10__12_), .D(_3748__bF_buf2), .Y(_4052_) );
NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_4050_), .B(_4051_), .C(_4052_), .Y(_4053_) );
NOR3X1 NOR3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_4045_), .B(_4049_), .C(_4053_), .Y(_4054_) );
AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf0), .B(_4032_), .C(_4041_), .D(_4054_), .Y(w_12_) );
XNOR2X1 XNOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__12_), .B(w_mem_inst_w_mem_13__12_), .Y(_4055_) );
XNOR2X1 XNOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__12_), .B(w_mem_inst_w_mem_2__12_), .Y(_4056_) );
XNOR2X1 XNOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_4055_), .B(_4056_), .Y(_4057_) );
INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__13_), .Y(_4058_) );
OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_3701_), .C(_3691__bF_buf4), .Y(_4059_) );
INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__13_), .Y(_4060_) );
NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__13_), .B(_3710__bF_buf4), .Y(_4061_) );
OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_4060_), .B(_3707_), .C(_4061_), .Y(_4062_) );
INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__13_), .Y(_4063_) );
INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__13_), .Y(_4064_) );
OAI22X1 OAI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(_4064_), .B(_3717__bF_buf2), .C(_4063_), .D(_3722__bF_buf2), .Y(_4065_) );
NOR3X1 NOR3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_4059_), .B(_4065_), .C(_4062_), .Y(_4066_) );
NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__13_), .B(_3727__bF_buf2), .Y(_4067_) );
NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__13_), .B(_3730__bF_buf2), .Y(_4068_) );
NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__13_), .B(_3732__bF_buf0), .Y(_4069_) );
NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_4068_), .B(_4069_), .C(_4067_), .Y(_4070_) );
AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf0), .B(w_mem_inst_w_mem_14__13_), .C(w_mem_inst_w_mem_7__13_), .D(_3736__bF_buf0), .Y(_4071_) );
NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__13_), .B(_3738__bF_buf4), .Y(_4072_) );
NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__13_), .B(_3740__bF_buf0), .Y(_4073_) );
NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_4072_), .B(_4073_), .C(_4071_), .Y(_4074_) );
NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__13_), .B(_3743_), .Y(_4075_) );
NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__13_), .B(_3745__bF_buf4), .Y(_4076_) );
AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf4), .B(w_mem_inst_w_mem_12__13_), .C(w_mem_inst_w_mem_10__13_), .D(_3748__bF_buf1), .Y(_4077_) );
NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_4075_), .B(_4076_), .C(_4077_), .Y(_4078_) );
NOR3X1 NOR3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_4070_), .B(_4074_), .C(_4078_), .Y(_4079_) );
AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf4), .B(_4057_), .C(_4066_), .D(_4079_), .Y(w_13_) );
XNOR2X1 XNOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__13_), .B(w_mem_inst_w_mem_13__13_), .Y(_4080_) );
XNOR2X1 XNOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__13_), .B(w_mem_inst_w_mem_2__13_), .Y(_4081_) );
XNOR2X1 XNOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_4080_), .B(_4081_), .Y(_4082_) );
INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__14_), .Y(_4083_) );
OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_4083_), .B(_3837_), .C(_3691__bF_buf3), .Y(_4084_) );
INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__14_), .Y(_4085_) );
INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__14_), .Y(_4086_) );
OAI22X1 OAI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_4086_), .B(_3838_), .C(_4085_), .D(_3763_), .Y(_4087_) );
INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__14_), .Y(_4088_) );
INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__14_), .Y(_4089_) );
OAI22X1 OAI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(_4088_), .B(_3717__bF_buf1), .C(_4089_), .D(_3756_), .Y(_4090_) );
NOR3X1 NOR3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_4084_), .B(_4090_), .C(_4087_), .Y(_4091_) );
NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__14_), .B(_3732__bF_buf4), .Y(_4092_) );
NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__14_), .B(_3730__bF_buf1), .Y(_4093_) );
NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__14_), .B(_3747__bF_buf3), .Y(_4094_) );
NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_4093_), .B(_4094_), .C(_4092_), .Y(_4095_) );
AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__14_), .B(_3710__bF_buf3), .C(w_mem_inst_w_mem_2__14_), .D(_3700__bF_buf3), .Y(_4096_) );
AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__14_), .B(_3745__bF_buf3), .C(w_mem_inst_w_mem_4__14_), .D(_3740__bF_buf3), .Y(_4097_) );
NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_4096_), .B(_4097_), .Y(_4098_) );
NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__14_), .B(_3706__bF_buf0), .Y(_4099_) );
NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__14_), .B(_3721_), .Y(_4100_) );
AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__14_), .B(_3738__bF_buf3), .C(w_mem_inst_w_mem_10__14_), .D(_3748__bF_buf0), .Y(_4101_) );
NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_4099_), .B(_4100_), .C(_4101_), .Y(_4102_) );
NOR3X1 NOR3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_4095_), .B(_4098_), .C(_4102_), .Y(_4103_) );
AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf3), .B(_4082_), .C(_4091_), .D(_4103_), .Y(w_14_) );
XNOR2X1 XNOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__14_), .B(w_mem_inst_w_mem_13__14_), .Y(_4104_) );
XNOR2X1 XNOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__14_), .B(w_mem_inst_w_mem_2__14_), .Y(_4105_) );
XNOR2X1 XNOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_4104_), .B(_4105_), .Y(_4106_) );
INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__15_), .Y(_4107_) );
OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_4107_), .B(_3833_), .C(_3691__bF_buf2), .Y(_4108_) );
INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__15_), .Y(_4109_) );
NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__15_), .B(_3747__bF_buf2), .Y(_4110_) );
OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_4109_), .B(_3717__bF_buf0), .C(_4110_), .Y(_4111_) );
INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__15_), .Y(_4112_) );
NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__15_), .B(_3710__bF_buf2), .Y(_4113_) );
OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_4112_), .B(_3707_), .C(_4113_), .Y(_4114_) );
NOR3X1 NOR3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_4111_), .B(_4108_), .C(_4114_), .Y(_4115_) );
NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__15_), .B(_3738__bF_buf2), .Y(_4116_) );
NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__15_), .B(_3730__bF_buf0), .Y(_4117_) );
NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__15_), .B(_3732__bF_buf3), .Y(_4118_) );
NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_4116_), .B(_4117_), .C(_4118_), .Y(_4119_) );
AOI22X1 AOI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__15_), .B(_3736__bF_buf3), .C(w_mem_inst_w_mem_8__15_), .D(_3721_), .Y(_4120_) );
NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__15_), .B(_3700__bF_buf2), .Y(_4121_) );
NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__15_), .B(_3748__bF_buf4), .Y(_4122_) );
NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_4121_), .B(_4122_), .C(_4120_), .Y(_4123_) );
AOI22X1 AOI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__15_), .B(_3745__bF_buf2), .C(w_mem_inst_w_mem_5__15_), .D(_3743_), .Y(_4124_) );
AOI22X1 AOI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__15_), .B(_3735__bF_buf4), .C(w_mem_inst_w_mem_9__15_), .D(_3727__bF_buf1), .Y(_4125_) );
NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_4124_), .B(_4125_), .Y(_4126_) );
NOR3X1 NOR3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_4119_), .B(_4126_), .C(_4123_), .Y(_4127_) );
AOI22X1 AOI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf2), .B(_4106_), .C(_4115_), .D(_4127_), .Y(w_15_) );
XNOR2X1 XNOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__15_), .B(w_mem_inst_w_mem_13__15_), .Y(_4128_) );
XNOR2X1 XNOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__15_), .B(w_mem_inst_w_mem_2__15_), .Y(_4129_) );
XNOR2X1 XNOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4128_), .B(_4129_), .Y(_4130_) );
INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__16_), .Y(_4131_) );
OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_4131_), .B(_3707_), .C(_3691__bF_buf1), .Y(_4132_) );
INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__16_), .Y(_4133_) );
INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__16_), .Y(_4134_) );
OAI22X1 OAI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(_4134_), .B(_3722__bF_buf1), .C(_4133_), .D(_3783_), .Y(_4135_) );
INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__16_), .Y(_4136_) );
INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__16_), .Y(_4137_) );
OAI22X1 OAI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_3838_), .C(_4137_), .D(_3764_), .Y(_4138_) );
NOR3X1 NOR3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_4138_), .B(_4132_), .C(_4135_), .Y(_4139_) );
NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__16_), .B(_3738__bF_buf1), .Y(_4140_) );
NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__16_), .B(_3745__bF_buf1), .Y(_4141_) );
NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__16_), .B(_3740__bF_buf2), .Y(_4142_) );
NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_4140_), .B(_4141_), .C(_4142_), .Y(_4143_) );
NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__16_), .B(_3727__bF_buf0), .Y(_4144_) );
NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__16_), .B(_3700__bF_buf1), .Y(_4145_) );
AOI22X1 AOI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__16_), .B(_3710__bF_buf1), .C(w_mem_inst_w_mem_1__16_), .D(_3732__bF_buf2), .Y(_4146_) );
NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_4144_), .B(_4145_), .C(_4146_), .Y(_4147_) );
AOI22X1 AOI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(w_mem_inst_w_mem_13__16_), .C(w_mem_inst_w_mem_14__16_), .D(_3735__bF_buf3), .Y(_4148_) );
NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__16_), .B(_3747__bF_buf1), .Y(_4149_) );
NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__16_), .B(_3743_), .Y(_4150_) );
NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_4149_), .B(_4150_), .C(_4148_), .Y(_4151_) );
NOR3X1 NOR3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_4143_), .B(_4151_), .C(_4147_), .Y(_4152_) );
AOI22X1 AOI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf1), .B(_4130_), .C(_4139_), .D(_4152_), .Y(w_16_) );
XNOR2X1 XNOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__16_), .B(w_mem_inst_w_mem_13__16_), .Y(_4153_) );
XNOR2X1 XNOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__16_), .B(w_mem_inst_w_mem_2__16_), .Y(_4154_) );
XNOR2X1 XNOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4153_), .B(_4154_), .Y(_4155_) );
INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__17_), .Y(_4156_) );
OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_4156_), .B(_3764_), .C(_3691__bF_buf0), .Y(_4157_) );
INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__17_), .Y(_4158_) );
INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__17_), .Y(_4159_) );
OAI22X1 OAI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(_4159_), .B(_3756_), .C(_4158_), .D(_3701_), .Y(_4160_) );
INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__17_), .Y(_4161_) );
INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__17_), .Y(_4162_) );
OAI22X1 OAI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_4162_), .B(_3717__bF_buf4), .C(_4161_), .D(_3722__bF_buf0), .Y(_4163_) );
NOR3X1 NOR3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_4157_), .B(_4160_), .C(_4163_), .Y(_4164_) );
NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__17_), .B(_3727__bF_buf3), .Y(_4165_) );
NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__17_), .B(_3732__bF_buf1), .Y(_4166_) );
NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__17_), .B(_3740__bF_buf1), .Y(_4167_) );
NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_4166_), .B(_4167_), .C(_4165_), .Y(_4168_) );
AOI22X1 AOI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf2), .B(w_mem_inst_w_mem_14__17_), .C(w_mem_inst_w_mem_7__17_), .D(_3736__bF_buf2), .Y(_4169_) );
NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__17_), .B(_3738__bF_buf0), .Y(_4170_) );
NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__17_), .B(_3706__bF_buf3), .Y(_4171_) );
NAND3X1 NAND3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_4170_), .B(_4171_), .C(_4169_), .Y(_4172_) );
AOI22X1 AOI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_3745__bF_buf0), .B(w_mem_inst_w_mem_11__17_), .C(w_mem_inst_w_mem_0__17_), .D(_3710__bF_buf0), .Y(_4173_) );
NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__17_), .B(_3747__bF_buf0), .Y(_4174_) );
NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__17_), .B(_3748__bF_buf3), .Y(_4175_) );
NAND3X1 NAND3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4174_), .B(_4175_), .C(_4173_), .Y(_4176_) );
NOR3X1 NOR3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_4168_), .B(_4172_), .C(_4176_), .Y(_4177_) );
AOI22X1 AOI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf0), .B(_4155_), .C(_4164_), .D(_4177_), .Y(w_17_) );
XNOR2X1 XNOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__17_), .B(w_mem_inst_w_mem_13__17_), .Y(_4178_) );
XNOR2X1 XNOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__17_), .B(w_mem_inst_w_mem_2__17_), .Y(_4179_) );
XNOR2X1 XNOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_4178_), .B(_4179_), .Y(_4180_) );
INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__18_), .Y(_4181_) );
OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_4181_), .B(_3701_), .C(_3691__bF_buf4), .Y(_4182_) );
INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__18_), .Y(_4183_) );
NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__18_), .B(_3710__bF_buf4), .Y(_4184_) );
OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_4183_), .B(_3756_), .C(_4184_), .Y(_4185_) );
INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__18_), .Y(_4186_) );
INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__18_), .Y(_4187_) );
OAI22X1 OAI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .B(_3717__bF_buf3), .C(_4186_), .D(_3722__bF_buf3), .Y(_4188_) );
NOR3X1 NOR3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_4185_), .B(_4182_), .C(_4188_), .Y(_4189_) );
NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__18_), .B(_3727__bF_buf2), .Y(_4190_) );
NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__18_), .B(_3730__bF_buf4), .Y(_4191_) );
NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__18_), .B(_3732__bF_buf0), .Y(_4192_) );
NAND3X1 NAND3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_4191_), .B(_4192_), .C(_4190_), .Y(_4193_) );
AOI22X1 AOI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf1), .B(w_mem_inst_w_mem_14__18_), .C(w_mem_inst_w_mem_7__18_), .D(_3736__bF_buf1), .Y(_4194_) );
NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__18_), .B(_3738__bF_buf4), .Y(_4195_) );
NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__18_), .B(_3740__bF_buf0), .Y(_4196_) );
NAND3X1 NAND3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_4195_), .B(_4196_), .C(_4194_), .Y(_4197_) );
NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__18_), .B(_3706__bF_buf2), .Y(_4198_) );
NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__18_), .B(_3745__bF_buf4), .Y(_4199_) );
AOI22X1 AOI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf4), .B(w_mem_inst_w_mem_12__18_), .C(w_mem_inst_w_mem_10__18_), .D(_3748__bF_buf2), .Y(_4200_) );
NAND3X1 NAND3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4198_), .B(_4199_), .C(_4200_), .Y(_4201_) );
NOR3X1 NOR3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_4193_), .B(_4197_), .C(_4201_), .Y(_4202_) );
AOI22X1 AOI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf4), .B(_4180_), .C(_4189_), .D(_4202_), .Y(w_18_) );
XNOR2X1 XNOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__18_), .B(w_mem_inst_w_mem_13__18_), .Y(_4203_) );
XNOR2X1 XNOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__18_), .B(w_mem_inst_w_mem_2__18_), .Y(_4204_) );
XNOR2X1 XNOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_4203_), .B(_4204_), .Y(_4205_) );
INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__19_), .Y(_4206_) );
OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_4206_), .B(_3833_), .C(_3691__bF_buf3), .Y(_4207_) );
INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__19_), .Y(_4208_) );
NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__19_), .B(_3710__bF_buf3), .Y(_4209_) );
OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_4208_), .B(_3707_), .C(_4209_), .Y(_4210_) );
INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__19_), .Y(_4211_) );
INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__19_), .Y(_4212_) );
OAI22X1 OAI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(_4212_), .B(_3717__bF_buf2), .C(_4211_), .D(_3722__bF_buf2), .Y(_4213_) );
NOR3X1 NOR3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_4207_), .B(_4213_), .C(_4210_), .Y(_4214_) );
NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__19_), .B(_3727__bF_buf1), .Y(_4215_) );
NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__19_), .B(_3730__bF_buf3), .Y(_4216_) );
NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__19_), .B(_3732__bF_buf4), .Y(_4217_) );
NAND3X1 NAND3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4216_), .B(_4217_), .C(_4215_), .Y(_4218_) );
AOI22X1 AOI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf0), .B(w_mem_inst_w_mem_14__19_), .C(w_mem_inst_w_mem_7__19_), .D(_3736__bF_buf0), .Y(_4219_) );
NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__19_), .B(_3738__bF_buf3), .Y(_4220_) );
NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__19_), .B(_3700__bF_buf0), .Y(_4221_) );
NAND3X1 NAND3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_4220_), .B(_4221_), .C(_4219_), .Y(_4222_) );
NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__19_), .B(_3743_), .Y(_4223_) );
NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__19_), .B(_3745__bF_buf3), .Y(_4224_) );
AOI22X1 AOI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf3), .B(w_mem_inst_w_mem_12__19_), .C(w_mem_inst_w_mem_10__19_), .D(_3748__bF_buf1), .Y(_4225_) );
NAND3X1 NAND3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_4223_), .B(_4224_), .C(_4225_), .Y(_4226_) );
NOR3X1 NOR3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_4218_), .B(_4222_), .C(_4226_), .Y(_4227_) );
AOI22X1 AOI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf3), .B(_4205_), .C(_4214_), .D(_4227_), .Y(w_19_) );
XNOR2X1 XNOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__19_), .B(w_mem_inst_w_mem_13__19_), .Y(_4228_) );
XNOR2X1 XNOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__19_), .B(w_mem_inst_w_mem_2__19_), .Y(_4229_) );
XNOR2X1 XNOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_4228_), .B(_4229_), .Y(_4230_) );
INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__20_), .Y(_4231_) );
OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_4231_), .B(_3833_), .C(_3691__bF_buf2), .Y(_4232_) );
INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__20_), .Y(_4233_) );
INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__20_), .Y(_4234_) );
OAI22X1 OAI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .B(_3838_), .C(_4233_), .D(_3763_), .Y(_4235_) );
INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__20_), .Y(_4236_) );
INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__20_), .Y(_4237_) );
OAI22X1 OAI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .B(_3717__bF_buf1), .C(_4237_), .D(_3756_), .Y(_4238_) );
NOR3X1 NOR3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_4238_), .B(_4232_), .C(_4235_), .Y(_4239_) );
NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__20_), .B(_3732__bF_buf3), .Y(_4240_) );
NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__20_), .B(_3730__bF_buf2), .Y(_4241_) );
NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__20_), .B(_3747__bF_buf2), .Y(_4242_) );
NAND3X1 NAND3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_4241_), .B(_4242_), .C(_4240_), .Y(_4243_) );
NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__20_), .B(_3710__bF_buf2), .Y(_4244_) );
NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__20_), .B(_3700__bF_buf3), .Y(_4245_) );
AOI22X1 AOI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf4), .B(w_mem_inst_w_mem_14__20_), .C(w_mem_inst_w_mem_11__20_), .D(_3745__bF_buf2), .Y(_4246_) );
NAND3X1 NAND3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_4244_), .B(_4245_), .C(_4246_), .Y(_4247_) );
NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__20_), .B(_3706__bF_buf1), .Y(_4248_) );
NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__20_), .B(_3721_), .Y(_4249_) );
AOI22X1 AOI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__20_), .B(_3738__bF_buf2), .C(w_mem_inst_w_mem_10__20_), .D(_3748__bF_buf0), .Y(_4250_) );
NAND3X1 NAND3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_4248_), .B(_4249_), .C(_4250_), .Y(_4251_) );
NOR3X1 NOR3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_4243_), .B(_4247_), .C(_4251_), .Y(_4252_) );
AOI22X1 AOI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf2), .B(_4230_), .C(_4239_), .D(_4252_), .Y(w_20_) );
XNOR2X1 XNOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__20_), .B(w_mem_inst_w_mem_13__20_), .Y(_4253_) );
XNOR2X1 XNOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__20_), .B(w_mem_inst_w_mem_2__20_), .Y(_4254_) );
XNOR2X1 XNOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_4253_), .B(_4254_), .Y(_4255_) );
INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__21_), .Y(_4256_) );
OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_4256_), .B(_3701_), .C(_3691__bF_buf1), .Y(_4257_) );
INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__21_), .Y(_4258_) );
NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__21_), .B(_3710__bF_buf1), .Y(_4259_) );
OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_4258_), .B(_3707_), .C(_4259_), .Y(_4260_) );
INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__21_), .Y(_4261_) );
INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__21_), .Y(_4262_) );
OAI22X1 OAI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_4262_), .B(_3717__bF_buf0), .C(_4261_), .D(_3722__bF_buf1), .Y(_4263_) );
NOR3X1 NOR3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_4257_), .B(_4263_), .C(_4260_), .Y(_4264_) );
NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__21_), .B(_3727__bF_buf0), .Y(_4265_) );
NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__21_), .B(_3730__bF_buf1), .Y(_4266_) );
NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__21_), .B(_3732__bF_buf2), .Y(_4267_) );
NAND3X1 NAND3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_4266_), .B(_4267_), .C(_4265_), .Y(_4268_) );
AOI22X1 AOI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf3), .B(w_mem_inst_w_mem_14__21_), .C(w_mem_inst_w_mem_7__21_), .D(_3736__bF_buf3), .Y(_4269_) );
NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__21_), .B(_3738__bF_buf1), .Y(_4270_) );
NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__21_), .B(_3740__bF_buf3), .Y(_4271_) );
NAND3X1 NAND3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_4270_), .B(_4271_), .C(_4269_), .Y(_4272_) );
NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__21_), .B(_3743_), .Y(_4273_) );
NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__21_), .B(_3745__bF_buf1), .Y(_4274_) );
AOI22X1 AOI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf1), .B(w_mem_inst_w_mem_12__21_), .C(w_mem_inst_w_mem_10__21_), .D(_3748__bF_buf4), .Y(_4275_) );
NAND3X1 NAND3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_4273_), .B(_4274_), .C(_4275_), .Y(_4276_) );
NOR3X1 NOR3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_4268_), .B(_4272_), .C(_4276_), .Y(_4277_) );
AOI22X1 AOI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf1), .B(_4255_), .C(_4264_), .D(_4277_), .Y(w_21_) );
XNOR2X1 XNOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__21_), .B(w_mem_inst_w_mem_13__21_), .Y(_4278_) );
XNOR2X1 XNOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__21_), .B(w_mem_inst_w_mem_2__21_), .Y(_4279_) );
XNOR2X1 XNOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_4278_), .B(_4279_), .Y(_4280_) );
INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__22_), .Y(_4281_) );
OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(_3837_), .C(_3691__bF_buf0), .Y(_4282_) );
INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__22_), .Y(_4283_) );
INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__22_), .Y(_4284_) );
OAI22X1 OAI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(_4284_), .B(_3838_), .C(_4283_), .D(_3763_), .Y(_4285_) );
INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__22_), .Y(_4286_) );
INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__22_), .Y(_4287_) );
OAI22X1 OAI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(_4286_), .B(_3717__bF_buf4), .C(_4287_), .D(_3756_), .Y(_4288_) );
NOR3X1 NOR3X1_39 ( .gnd(gnd), .vdd(vdd), .A(_4282_), .B(_4288_), .C(_4285_), .Y(_4289_) );
NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__22_), .B(_3732__bF_buf1), .Y(_4290_) );
NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__22_), .B(_3730__bF_buf0), .Y(_4291_) );
NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__22_), .B(_3747__bF_buf0), .Y(_4292_) );
NAND3X1 NAND3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_4291_), .B(_4292_), .C(_4290_), .Y(_4293_) );
AOI22X1 AOI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__22_), .B(_3710__bF_buf0), .C(w_mem_inst_w_mem_2__22_), .D(_3700__bF_buf2), .Y(_4294_) );
AOI22X1 AOI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__22_), .B(_3745__bF_buf0), .C(w_mem_inst_w_mem_4__22_), .D(_3740__bF_buf2), .Y(_4295_) );
NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_4294_), .B(_4295_), .Y(_4296_) );
NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__22_), .B(_3706__bF_buf0), .Y(_4297_) );
NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__22_), .B(_3721_), .Y(_4298_) );
AOI22X1 AOI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__22_), .B(_3738__bF_buf0), .C(w_mem_inst_w_mem_10__22_), .D(_3748__bF_buf3), .Y(_4299_) );
NAND3X1 NAND3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_4297_), .B(_4298_), .C(_4299_), .Y(_4300_) );
NOR3X1 NOR3X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4293_), .B(_4296_), .C(_4300_), .Y(_4301_) );
AOI22X1 AOI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf0), .B(_4280_), .C(_4289_), .D(_4301_), .Y(w_22_) );
XNOR2X1 XNOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__22_), .B(w_mem_inst_w_mem_13__22_), .Y(_4302_) );
XNOR2X1 XNOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__22_), .B(w_mem_inst_w_mem_2__22_), .Y(_4303_) );
XNOR2X1 XNOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_4302_), .B(_4303_), .Y(_4304_) );
INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__23_), .Y(_4305_) );
OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_4305_), .B(_3833_), .C(_3691__bF_buf4), .Y(_4306_) );
INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__23_), .Y(_4307_) );
NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__23_), .B(_3747__bF_buf4), .Y(_4308_) );
OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_4307_), .B(_3717__bF_buf3), .C(_4308_), .Y(_4309_) );
INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__23_), .Y(_4310_) );
NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__23_), .B(_3710__bF_buf4), .Y(_4311_) );
OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_4310_), .B(_3707_), .C(_4311_), .Y(_4312_) );
NOR3X1 NOR3X1_41 ( .gnd(gnd), .vdd(vdd), .A(_4309_), .B(_4306_), .C(_4312_), .Y(_4313_) );
NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__23_), .B(_3738__bF_buf4), .Y(_4314_) );
NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__23_), .B(_3730__bF_buf4), .Y(_4315_) );
NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__23_), .B(_3732__bF_buf0), .Y(_4316_) );
NAND3X1 NAND3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_4314_), .B(_4315_), .C(_4316_), .Y(_4317_) );
AOI22X1 AOI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__23_), .B(_3736__bF_buf2), .C(w_mem_inst_w_mem_8__23_), .D(_3721_), .Y(_4318_) );
NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__23_), .B(_3700__bF_buf1), .Y(_4319_) );
NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__23_), .B(_3748__bF_buf2), .Y(_4320_) );
NAND3X1 NAND3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_4319_), .B(_4320_), .C(_4318_), .Y(_4321_) );
AOI22X1 AOI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__23_), .B(_3745__bF_buf4), .C(w_mem_inst_w_mem_5__23_), .D(_3743_), .Y(_4322_) );
AOI22X1 AOI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__23_), .B(_3735__bF_buf2), .C(w_mem_inst_w_mem_9__23_), .D(_3727__bF_buf3), .Y(_4323_) );
NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_4322_), .B(_4323_), .Y(_4324_) );
NOR3X1 NOR3X1_42 ( .gnd(gnd), .vdd(vdd), .A(_4317_), .B(_4324_), .C(_4321_), .Y(_4325_) );
AOI22X1 AOI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf4), .B(_4304_), .C(_4313_), .D(_4325_), .Y(w_23_) );
XNOR2X1 XNOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__23_), .B(w_mem_inst_w_mem_13__23_), .Y(_4326_) );
XNOR2X1 XNOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__23_), .B(w_mem_inst_w_mem_2__23_), .Y(_4327_) );
XNOR2X1 XNOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_4326_), .B(_4327_), .Y(_4328_) );
INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__24_), .Y(_4329_) );
OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_4329_), .B(_3707_), .C(_3691__bF_buf3), .Y(_4330_) );
INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__24_), .Y(_4331_) );
INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__24_), .Y(_4332_) );
OAI22X1 OAI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .B(_3722__bF_buf0), .C(_4331_), .D(_3783_), .Y(_4333_) );
INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__24_), .Y(_4334_) );
INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__24_), .Y(_4335_) );
OAI22X1 OAI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(_4334_), .B(_3838_), .C(_4335_), .D(_3764_), .Y(_4336_) );
NOR3X1 NOR3X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4336_), .B(_4330_), .C(_4333_), .Y(_4337_) );
NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__24_), .B(_3738__bF_buf3), .Y(_4338_) );
NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__24_), .B(_3745__bF_buf3), .Y(_4339_) );
NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__24_), .B(_3740__bF_buf1), .Y(_4340_) );
NAND3X1 NAND3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_4338_), .B(_4339_), .C(_4340_), .Y(_4341_) );
NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__24_), .B(_3727__bF_buf2), .Y(_4342_) );
NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__24_), .B(_3700__bF_buf0), .Y(_4343_) );
AOI22X1 AOI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__24_), .B(_3710__bF_buf3), .C(w_mem_inst_w_mem_1__24_), .D(_3732__bF_buf4), .Y(_4344_) );
NAND3X1 NAND3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_4342_), .B(_4343_), .C(_4344_), .Y(_4345_) );
AOI22X1 AOI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(w_mem_inst_w_mem_13__24_), .C(w_mem_inst_w_mem_14__24_), .D(_3735__bF_buf1), .Y(_4346_) );
NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__24_), .B(_3747__bF_buf3), .Y(_4347_) );
NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__24_), .B(_3743_), .Y(_4348_) );
NAND3X1 NAND3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_4347_), .B(_4348_), .C(_4346_), .Y(_4349_) );
NOR3X1 NOR3X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4341_), .B(_4349_), .C(_4345_), .Y(_4350_) );
AOI22X1 AOI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf3), .B(_4328_), .C(_4337_), .D(_4350_), .Y(w_24_) );
XNOR2X1 XNOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__24_), .B(w_mem_inst_w_mem_13__24_), .Y(_4351_) );
XNOR2X1 XNOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__24_), .B(w_mem_inst_w_mem_2__24_), .Y(_4352_) );
XNOR2X1 XNOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_4351_), .B(_4352_), .Y(_4353_) );
INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__25_), .Y(_4354_) );
OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .B(_3764_), .C(_3691__bF_buf2), .Y(_4355_) );
INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__25_), .Y(_4356_) );
INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__25_), .Y(_4357_) );
OAI22X1 OAI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_4357_), .B(_3756_), .C(_4356_), .D(_3701_), .Y(_4358_) );
INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__25_), .Y(_4359_) );
INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__25_), .Y(_4360_) );
OAI22X1 OAI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(_4360_), .B(_3717__bF_buf2), .C(_4359_), .D(_3722__bF_buf3), .Y(_4361_) );
NOR3X1 NOR3X1_45 ( .gnd(gnd), .vdd(vdd), .A(_4355_), .B(_4358_), .C(_4361_), .Y(_4362_) );
NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__25_), .B(_3727__bF_buf1), .Y(_4363_) );
NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__25_), .B(_3732__bF_buf3), .Y(_4364_) );
NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__25_), .B(_3740__bF_buf0), .Y(_4365_) );
NAND3X1 NAND3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_4364_), .B(_4365_), .C(_4363_), .Y(_4366_) );
AOI22X1 AOI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf0), .B(w_mem_inst_w_mem_14__25_), .C(w_mem_inst_w_mem_7__25_), .D(_3736__bF_buf1), .Y(_4367_) );
NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__25_), .B(_3738__bF_buf2), .Y(_4368_) );
NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__25_), .B(_3706__bF_buf3), .Y(_4369_) );
NAND3X1 NAND3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_4368_), .B(_4369_), .C(_4367_), .Y(_4370_) );
AOI22X1 AOI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_3745__bF_buf2), .B(w_mem_inst_w_mem_11__25_), .C(w_mem_inst_w_mem_0__25_), .D(_3710__bF_buf2), .Y(_4371_) );
NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__25_), .B(_3747__bF_buf2), .Y(_4372_) );
NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__25_), .B(_3748__bF_buf1), .Y(_4373_) );
NAND3X1 NAND3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_4372_), .B(_4373_), .C(_4371_), .Y(_4374_) );
NOR3X1 NOR3X1_46 ( .gnd(gnd), .vdd(vdd), .A(_4366_), .B(_4370_), .C(_4374_), .Y(_4375_) );
AOI22X1 AOI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf2), .B(_4353_), .C(_4362_), .D(_4375_), .Y(w_25_) );
XNOR2X1 XNOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__25_), .B(w_mem_inst_w_mem_13__25_), .Y(_4376_) );
XNOR2X1 XNOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__25_), .B(w_mem_inst_w_mem_2__25_), .Y(_4377_) );
XNOR2X1 XNOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_4376_), .B(_4377_), .Y(_4378_) );
INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__26_), .Y(_4379_) );
OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_4379_), .B(_3701_), .C(_3691__bF_buf1), .Y(_4380_) );
INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__26_), .Y(_4381_) );
NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__26_), .B(_3710__bF_buf1), .Y(_4382_) );
OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4381_), .B(_3756_), .C(_4382_), .Y(_4383_) );
INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__26_), .Y(_4384_) );
INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__26_), .Y(_4385_) );
OAI22X1 OAI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(_4385_), .B(_3717__bF_buf1), .C(_4384_), .D(_3722__bF_buf2), .Y(_4386_) );
NOR3X1 NOR3X1_47 ( .gnd(gnd), .vdd(vdd), .A(_4383_), .B(_4380_), .C(_4386_), .Y(_4387_) );
NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__26_), .B(_3727__bF_buf0), .Y(_4388_) );
NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__26_), .B(_3730__bF_buf3), .Y(_4389_) );
NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__26_), .B(_3732__bF_buf2), .Y(_4390_) );
NAND3X1 NAND3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_4389_), .B(_4390_), .C(_4388_), .Y(_4391_) );
AOI22X1 AOI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf4), .B(w_mem_inst_w_mem_14__26_), .C(w_mem_inst_w_mem_7__26_), .D(_3736__bF_buf0), .Y(_4392_) );
NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__26_), .B(_3738__bF_buf1), .Y(_4393_) );
NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__26_), .B(_3740__bF_buf3), .Y(_4394_) );
NAND3X1 NAND3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_4393_), .B(_4394_), .C(_4392_), .Y(_4395_) );
NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__26_), .B(_3706__bF_buf2), .Y(_4396_) );
NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__26_), .B(_3745__bF_buf1), .Y(_4397_) );
AOI22X1 AOI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf1), .B(w_mem_inst_w_mem_12__26_), .C(w_mem_inst_w_mem_10__26_), .D(_3748__bF_buf0), .Y(_4398_) );
NAND3X1 NAND3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_4396_), .B(_4397_), .C(_4398_), .Y(_4399_) );
NOR3X1 NOR3X1_48 ( .gnd(gnd), .vdd(vdd), .A(_4391_), .B(_4395_), .C(_4399_), .Y(_4400_) );
AOI22X1 AOI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf1), .B(_4378_), .C(_4387_), .D(_4400_), .Y(w_26_) );
XNOR2X1 XNOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__26_), .B(w_mem_inst_w_mem_13__26_), .Y(_4401_) );
XNOR2X1 XNOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__26_), .B(w_mem_inst_w_mem_2__26_), .Y(_4402_) );
XNOR2X1 XNOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_4401_), .B(_4402_), .Y(_4403_) );
INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__27_), .Y(_4404_) );
OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_4404_), .B(_3833_), .C(_3691__bF_buf0), .Y(_4405_) );
INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__27_), .Y(_4406_) );
NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__27_), .B(_3710__bF_buf0), .Y(_4407_) );
OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_4406_), .B(_3707_), .C(_4407_), .Y(_4408_) );
INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__27_), .Y(_4409_) );
INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__27_), .Y(_4410_) );
OAI22X1 OAI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_4410_), .B(_3717__bF_buf0), .C(_4409_), .D(_3722__bF_buf1), .Y(_4411_) );
NOR3X1 NOR3X1_49 ( .gnd(gnd), .vdd(vdd), .A(_4405_), .B(_4411_), .C(_4408_), .Y(_4412_) );
NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__27_), .B(_3727__bF_buf3), .Y(_4413_) );
NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__27_), .B(_3730__bF_buf2), .Y(_4414_) );
NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__27_), .B(_3732__bF_buf1), .Y(_4415_) );
NAND3X1 NAND3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_4414_), .B(_4415_), .C(_4413_), .Y(_4416_) );
AOI22X1 AOI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf3), .B(w_mem_inst_w_mem_14__27_), .C(w_mem_inst_w_mem_7__27_), .D(_3736__bF_buf3), .Y(_4417_) );
NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__27_), .B(_3738__bF_buf0), .Y(_4418_) );
NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__27_), .B(_3700__bF_buf3), .Y(_4419_) );
NAND3X1 NAND3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_4418_), .B(_4419_), .C(_4417_), .Y(_4420_) );
NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__27_), .B(_3743_), .Y(_4421_) );
NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__27_), .B(_3745__bF_buf0), .Y(_4422_) );
AOI22X1 AOI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf0), .B(w_mem_inst_w_mem_12__27_), .C(w_mem_inst_w_mem_10__27_), .D(_3748__bF_buf4), .Y(_4423_) );
NAND3X1 NAND3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_4421_), .B(_4422_), .C(_4423_), .Y(_4424_) );
NOR3X1 NOR3X1_50 ( .gnd(gnd), .vdd(vdd), .A(_4416_), .B(_4420_), .C(_4424_), .Y(_4425_) );
AOI22X1 AOI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf0), .B(_4403_), .C(_4412_), .D(_4425_), .Y(w_27_) );
XNOR2X1 XNOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__27_), .B(w_mem_inst_w_mem_13__27_), .Y(_4426_) );
XNOR2X1 XNOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__27_), .B(w_mem_inst_w_mem_2__27_), .Y(_4427_) );
XNOR2X1 XNOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_4426_), .B(_4427_), .Y(_4428_) );
INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__28_), .Y(_4429_) );
OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_3833_), .C(_3691__bF_buf4), .Y(_4430_) );
INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__28_), .Y(_4431_) );
INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__28_), .Y(_4432_) );
OAI22X1 OAI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(_4432_), .B(_3838_), .C(_4431_), .D(_3763_), .Y(_4433_) );
INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__28_), .Y(_4434_) );
INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__28_), .Y(_4435_) );
OAI22X1 OAI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_3717__bF_buf4), .C(_4435_), .D(_3756_), .Y(_4436_) );
NOR3X1 NOR3X1_51 ( .gnd(gnd), .vdd(vdd), .A(_4436_), .B(_4430_), .C(_4433_), .Y(_4437_) );
NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__28_), .B(_3732__bF_buf0), .Y(_4438_) );
NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__28_), .B(_3730__bF_buf1), .Y(_4439_) );
NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__28_), .B(_3747__bF_buf4), .Y(_4440_) );
NAND3X1 NAND3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_4439_), .B(_4440_), .C(_4438_), .Y(_4441_) );
NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__28_), .B(_3710__bF_buf4), .Y(_4442_) );
NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__28_), .B(_3700__bF_buf2), .Y(_4443_) );
AOI22X1 AOI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf2), .B(w_mem_inst_w_mem_14__28_), .C(w_mem_inst_w_mem_11__28_), .D(_3745__bF_buf4), .Y(_4444_) );
NAND3X1 NAND3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_4442_), .B(_4443_), .C(_4444_), .Y(_4445_) );
NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__28_), .B(_3706__bF_buf1), .Y(_4446_) );
NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__28_), .B(_3721_), .Y(_4447_) );
AOI22X1 AOI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__28_), .B(_3738__bF_buf4), .C(w_mem_inst_w_mem_10__28_), .D(_3748__bF_buf3), .Y(_4448_) );
NAND3X1 NAND3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_4446_), .B(_4447_), .C(_4448_), .Y(_4449_) );
NOR3X1 NOR3X1_52 ( .gnd(gnd), .vdd(vdd), .A(_4441_), .B(_4445_), .C(_4449_), .Y(_4450_) );
AOI22X1 AOI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf4), .B(_4428_), .C(_4437_), .D(_4450_), .Y(w_28_) );
XNOR2X1 XNOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__28_), .B(w_mem_inst_w_mem_13__28_), .Y(_4451_) );
XNOR2X1 XNOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__28_), .B(w_mem_inst_w_mem_2__28_), .Y(_4452_) );
XNOR2X1 XNOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_4451_), .B(_4452_), .Y(_4453_) );
INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__29_), .Y(_4454_) );
OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_4454_), .B(_3701_), .C(_3691__bF_buf3), .Y(_4455_) );
INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__29_), .Y(_4456_) );
NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__29_), .B(_3710__bF_buf3), .Y(_4457_) );
OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_4456_), .B(_3707_), .C(_4457_), .Y(_4458_) );
INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__29_), .Y(_4459_) );
INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__29_), .Y(_4460_) );
OAI22X1 OAI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(_4460_), .B(_3717__bF_buf3), .C(_4459_), .D(_3722__bF_buf0), .Y(_4461_) );
NOR3X1 NOR3X1_53 ( .gnd(gnd), .vdd(vdd), .A(_4455_), .B(_4461_), .C(_4458_), .Y(_4462_) );
NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__29_), .B(_3727__bF_buf2), .Y(_4463_) );
NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__29_), .B(_3730__bF_buf0), .Y(_4464_) );
NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__29_), .B(_3732__bF_buf4), .Y(_4465_) );
NAND3X1 NAND3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_4464_), .B(_4465_), .C(_4463_), .Y(_4466_) );
AOI22X1 AOI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf1), .B(w_mem_inst_w_mem_14__29_), .C(w_mem_inst_w_mem_7__29_), .D(_3736__bF_buf2), .Y(_4467_) );
NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__29_), .B(_3738__bF_buf3), .Y(_4468_) );
NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__29_), .B(_3740__bF_buf2), .Y(_4469_) );
NAND3X1 NAND3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_4468_), .B(_4469_), .C(_4467_), .Y(_4470_) );
NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__29_), .B(_3743_), .Y(_4471_) );
NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__29_), .B(_3745__bF_buf3), .Y(_4472_) );
AOI22X1 AOI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf3), .B(w_mem_inst_w_mem_12__29_), .C(w_mem_inst_w_mem_10__29_), .D(_3748__bF_buf2), .Y(_4473_) );
NAND3X1 NAND3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_4471_), .B(_4472_), .C(_4473_), .Y(_4474_) );
NOR3X1 NOR3X1_54 ( .gnd(gnd), .vdd(vdd), .A(_4466_), .B(_4470_), .C(_4474_), .Y(_4475_) );
AOI22X1 AOI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf3), .B(_4453_), .C(_4462_), .D(_4475_), .Y(w_29_) );
XNOR2X1 XNOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__29_), .B(w_mem_inst_w_mem_13__29_), .Y(_4476_) );
XNOR2X1 XNOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__29_), .B(w_mem_inst_w_mem_2__29_), .Y(_4477_) );
XNOR2X1 XNOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_4476_), .B(_4477_), .Y(_4478_) );
INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__30_), .Y(_4479_) );
OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_3837_), .C(_3691__bF_buf2), .Y(_4480_) );
INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__30_), .Y(_4481_) );
INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__30_), .Y(_4482_) );
OAI22X1 OAI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_3838_), .C(_4481_), .D(_3763_), .Y(_4483_) );
INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__30_), .Y(_4484_) );
INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__30_), .Y(_4485_) );
OAI22X1 OAI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_4484_), .B(_3717__bF_buf2), .C(_4485_), .D(_3756_), .Y(_4486_) );
NOR3X1 NOR3X1_55 ( .gnd(gnd), .vdd(vdd), .A(_4480_), .B(_4486_), .C(_4483_), .Y(_4487_) );
NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__30_), .B(_3732__bF_buf3), .Y(_4488_) );
NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__30_), .B(_3730__bF_buf4), .Y(_4489_) );
NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__30_), .B(_3747__bF_buf2), .Y(_4490_) );
NAND3X1 NAND3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_4489_), .B(_4490_), .C(_4488_), .Y(_4491_) );
AOI22X1 AOI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__30_), .B(_3710__bF_buf2), .C(w_mem_inst_w_mem_2__30_), .D(_3700__bF_buf1), .Y(_4492_) );
AOI22X1 AOI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__30_), .B(_3745__bF_buf2), .C(w_mem_inst_w_mem_4__30_), .D(_3740__bF_buf1), .Y(_4493_) );
NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_4492_), .B(_4493_), .Y(_4494_) );
NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__30_), .B(_3706__bF_buf0), .Y(_4495_) );
NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__30_), .B(_3721_), .Y(_4496_) );
AOI22X1 AOI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__30_), .B(_3738__bF_buf2), .C(w_mem_inst_w_mem_10__30_), .D(_3748__bF_buf1), .Y(_4497_) );
NAND3X1 NAND3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_4495_), .B(_4496_), .C(_4497_), .Y(_4498_) );
NOR3X1 NOR3X1_56 ( .gnd(gnd), .vdd(vdd), .A(_4491_), .B(_4494_), .C(_4498_), .Y(_4499_) );
AOI22X1 AOI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf2), .B(_4478_), .C(_4487_), .D(_4499_), .Y(w_30_) );
XNOR2X1 XNOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__30_), .B(w_mem_inst_w_mem_13__30_), .Y(_4500_) );
XNOR2X1 XNOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__30_), .B(w_mem_inst_w_mem_2__30_), .Y(_4501_) );
XNOR2X1 XNOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_4500_), .B(_4501_), .Y(_4502_) );
INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__31_), .Y(_4503_) );
OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_4503_), .B(_3833_), .C(_3691__bF_buf1), .Y(_4504_) );
INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__31_), .Y(_4505_) );
INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__31_), .Y(_4506_) );
OAI22X1 OAI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_3838_), .C(_4506_), .D(_3837_), .Y(_4507_) );
INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__31_), .Y(_4508_) );
INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__31_), .Y(_4509_) );
OAI22X1 OAI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_4508_), .B(_3763_), .C(_4509_), .D(_3707_), .Y(_4510_) );
NOR3X1 NOR3X1_57 ( .gnd(gnd), .vdd(vdd), .A(_4507_), .B(_4504_), .C(_4510_), .Y(_4511_) );
NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__31_), .B(_3732__bF_buf2), .Y(_4512_) );
NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__31_), .B(_3730__bF_buf3), .Y(_4513_) );
NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__31_), .B(_3748__bF_buf0), .Y(_4514_) );
NAND3X1 NAND3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_4513_), .B(_4512_), .C(_4514_), .Y(_4515_) );
AOI22X1 AOI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__31_), .B(_3710__bF_buf1), .C(w_mem_inst_w_mem_2__31_), .D(_3700__bF_buf0), .Y(_4516_) );
NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__31_), .B(_3745__bF_buf1), .Y(_4517_) );
NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__31_), .B(_3721_), .Y(_4518_) );
NAND3X1 NAND3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_4517_), .B(_4518_), .C(_4516_), .Y(_4519_) );
NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__31_), .B(_3743_), .Y(_4520_) );
NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__31_), .B(_3747__bF_buf1), .Y(_4521_) );
AOI22X1 AOI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__31_), .B(_3738__bF_buf1), .C(w_mem_inst_w_mem_13__31_), .D(_3716_), .Y(_4522_) );
NAND3X1 NAND3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_4521_), .B(_4522_), .C(_4520_), .Y(_4523_) );
NOR3X1 NOR3X1_58 ( .gnd(gnd), .vdd(vdd), .A(_4515_), .B(_4523_), .C(_4519_), .Y(_4524_) );
AOI22X1 AOI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf1), .B(_4502_), .C(_4511_), .D(_4524_), .Y(w_31_) );
INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .Y(_4525_) );
AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(w_mem_inst_sha1_w_mem_ctrl_reg), .Y(_4526_) );
INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(_4526_), .Y(_4527_) );
OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_sha1_w_mem_ctrl_reg), .B(_4525_), .C(_4527_), .Y(_4528_) );
NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_3698_), .B(_4526_), .Y(_4529_) );
OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_3698_), .B(_4528_), .C(_4529_), .Y(_3671__0_) );
NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3726_), .Y(_4530_) );
NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_4526_), .B(_4530_), .Y(_4531_) );
OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(_4528_), .C(_4531_), .Y(_3671__1_) );
INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(_3729_), .Y(_4532_) );
NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_2_), .B(_4532_), .Y(_4533_) );
OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_3725_), .B(_3698_), .C(_3719_), .Y(_4534_) );
NAND3X1 NAND3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_4526_), .B(_4534_), .C(_4533_), .Y(_4535_) );
OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_3719_), .B(_4528_), .C(_4535_), .Y(_3671__2_) );
AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_4533_), .B(w_mem_inst_w_ctr_reg_3_), .C(_3736__bF_buf1), .Y(_4536_) );
OAI22X1 OAI22X1_41 ( .gnd(gnd), .vdd(vdd), .A(_3704_), .B(_4528_), .C(_4527_), .D(_4536_), .Y(_3671__3_) );
OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_sha1_w_mem_ctrl_reg), .B(_4525_), .C(w_mem_inst_w_ctr_reg_4_), .Y(_4537_) );
NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_4526_), .B(_3738__bF_buf0), .Y(_4538_) );
NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_3688_), .B(_4538_), .Y(_4539_) );
AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_4537_), .B(_4538_), .C(_4539_), .Y(_3671__4_) );
OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_sha1_w_mem_ctrl_reg), .B(_4525_), .C(w_mem_inst_w_ctr_reg_5_), .Y(_4540_) );
MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_5_), .B(_4540_), .S(_4539_), .Y(_3671__5_) );
NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_5_), .B(_4539_), .Y(_4541_) );
OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_sha1_w_mem_ctrl_reg), .B(_4525_), .C(w_mem_inst_w_ctr_reg_6_), .Y(_4542_) );
MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_4542_), .B(w_mem_inst_w_ctr_reg_6_), .S(_4541_), .Y(_3671__6_) );
INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(_3738__bF_buf4), .Y(_4543_) );
NAND3X1 NAND3X1_81 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_6_), .B(_3688_), .C(_3689_), .Y(_4544_) );
OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_4544_), .B(_4543_), .C(w_mem_inst_sha1_w_mem_ctrl_reg), .Y(_4545_) );
OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_sha1_w_mem_ctrl_reg), .B(_4525_), .C(_4545_), .Y(_3670_) );
INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__0_), .Y(_4546_) );
OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_6_), .B(_3690_), .C(_4525_), .Y(_4547_) );
NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(_3692__bF_buf0), .Y(_4548_) );
AOI22X1 AOI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[480]), .C(w_mem_inst_w_mem_0__0_), .D(_4548__bF_buf63), .Y(_4549_) );
OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_4546_), .B(_4547__bF_buf63), .C(_4549_), .Y(_3672__0_) );
INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__1_), .Y(_4550_) );
AOI22X1 AOI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[481]), .C(w_mem_inst_w_mem_0__1_), .D(_4548__bF_buf62), .Y(_4551_) );
OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_4550_), .B(_4547__bF_buf62), .C(_4551_), .Y(_3672__1_) );
AOI22X1 AOI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[482]), .C(w_mem_inst_w_mem_0__2_), .D(_4548__bF_buf61), .Y(_4552_) );
OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3788_), .B(_4547__bF_buf61), .C(_4552_), .Y(_3672__2_) );
INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__3_), .Y(_4553_) );
AOI22X1 AOI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[483]), .C(w_mem_inst_w_mem_0__3_), .D(_4548__bF_buf60), .Y(_4554_) );
OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_4553_), .B(_4547__bF_buf60), .C(_4554_), .Y(_3672__3_) );
INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__4_), .Y(_4555_) );
AOI22X1 AOI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[484]), .C(w_mem_inst_w_mem_0__4_), .D(_4548__bF_buf59), .Y(_4556_) );
OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_4555_), .B(_4547__bF_buf59), .C(_4556_), .Y(_3672__4_) );
AOI22X1 AOI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[485]), .C(w_mem_inst_w_mem_0__5_), .D(_4548__bF_buf58), .Y(_4557_) );
OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_3865_), .B(_4547__bF_buf58), .C(_4557_), .Y(_3672__5_) );
INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__6_), .Y(_4558_) );
AOI22X1 AOI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[486]), .C(w_mem_inst_w_mem_0__6_), .D(_4548__bF_buf57), .Y(_4559_) );
OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_4558_), .B(_4547__bF_buf57), .C(_4559_), .Y(_3672__6_) );
INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__7_), .Y(_4560_) );
AOI22X1 AOI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[487]), .C(w_mem_inst_w_mem_0__7_), .D(_4548__bF_buf56), .Y(_4561_) );
OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_4560_), .B(_4547__bF_buf56), .C(_4561_), .Y(_3672__7_) );
INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__8_), .Y(_4562_) );
AOI22X1 AOI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[488]), .C(w_mem_inst_w_mem_0__8_), .D(_4548__bF_buf55), .Y(_4563_) );
OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_4562_), .B(_4547__bF_buf55), .C(_4563_), .Y(_3672__8_) );
INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__9_), .Y(_4564_) );
AOI22X1 AOI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[489]), .C(w_mem_inst_w_mem_0__9_), .D(_4548__bF_buf54), .Y(_4565_) );
OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_4564_), .B(_4547__bF_buf54), .C(_4565_), .Y(_3672__9_) );
INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__10_), .Y(_4566_) );
AOI22X1 AOI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[490]), .C(w_mem_inst_w_mem_0__10_), .D(_4548__bF_buf53), .Y(_4567_) );
OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_4566_), .B(_4547__bF_buf53), .C(_4567_), .Y(_3672__10_) );
INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__11_), .Y(_4568_) );
AOI22X1 AOI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[491]), .C(w_mem_inst_w_mem_0__11_), .D(_4548__bF_buf52), .Y(_4569_) );
OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_4568_), .B(_4547__bF_buf52), .C(_4569_), .Y(_3672__11_) );
INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__12_), .Y(_4570_) );
AOI22X1 AOI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[492]), .C(w_mem_inst_w_mem_0__12_), .D(_4548__bF_buf51), .Y(_4571_) );
OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_4570_), .B(_4547__bF_buf51), .C(_4571_), .Y(_3672__12_) );
INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__13_), .Y(_4572_) );
AOI22X1 AOI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[493]), .C(w_mem_inst_w_mem_0__13_), .D(_4548__bF_buf50), .Y(_4573_) );
OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_4572_), .B(_4547__bF_buf50), .C(_4573_), .Y(_3672__13_) );
INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__14_), .Y(_4574_) );
AOI22X1 AOI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[494]), .C(w_mem_inst_w_mem_0__14_), .D(_4548__bF_buf49), .Y(_4575_) );
OAI21X1 OAI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_4574_), .B(_4547__bF_buf49), .C(_4575_), .Y(_3672__14_) );
INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__15_), .Y(_4576_) );
AOI22X1 AOI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[495]), .C(w_mem_inst_w_mem_0__15_), .D(_4548__bF_buf48), .Y(_4577_) );
OAI21X1 OAI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_4576_), .B(_4547__bF_buf48), .C(_4577_), .Y(_3672__15_) );
INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__16_), .Y(_4578_) );
AOI22X1 AOI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[496]), .C(w_mem_inst_w_mem_0__16_), .D(_4548__bF_buf47), .Y(_4579_) );
OAI21X1 OAI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_4578_), .B(_4547__bF_buf47), .C(_4579_), .Y(_3672__16_) );
INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__17_), .Y(_4580_) );
AOI22X1 AOI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[497]), .C(w_mem_inst_w_mem_0__17_), .D(_4548__bF_buf46), .Y(_4581_) );
OAI21X1 OAI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_4580_), .B(_4547__bF_buf46), .C(_4581_), .Y(_3672__17_) );
INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__18_), .Y(_4582_) );
AOI22X1 AOI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[498]), .C(w_mem_inst_w_mem_0__18_), .D(_4548__bF_buf45), .Y(_4583_) );
OAI21X1 OAI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_4582_), .B(_4547__bF_buf45), .C(_4583_), .Y(_3672__18_) );
INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__19_), .Y(_4584_) );
AOI22X1 AOI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[499]), .C(w_mem_inst_w_mem_0__19_), .D(_4548__bF_buf44), .Y(_4585_) );
OAI21X1 OAI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_4584_), .B(_4547__bF_buf44), .C(_4585_), .Y(_3672__19_) );
INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__20_), .Y(_4586_) );
AOI22X1 AOI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[500]), .C(w_mem_inst_w_mem_0__20_), .D(_4548__bF_buf43), .Y(_4587_) );
OAI21X1 OAI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_4586_), .B(_4547__bF_buf43), .C(_4587_), .Y(_3672__20_) );
INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__21_), .Y(_4588_) );
AOI22X1 AOI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[501]), .C(w_mem_inst_w_mem_0__21_), .D(_4548__bF_buf42), .Y(_4589_) );
OAI21X1 OAI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_4588_), .B(_4547__bF_buf42), .C(_4589_), .Y(_3672__21_) );
INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__22_), .Y(_4590_) );
AOI22X1 AOI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[502]), .C(w_mem_inst_w_mem_0__22_), .D(_4548__bF_buf41), .Y(_4591_) );
OAI21X1 OAI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_4590_), .B(_4547__bF_buf41), .C(_4591_), .Y(_3672__22_) );
INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__23_), .Y(_4592_) );
AOI22X1 AOI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[503]), .C(w_mem_inst_w_mem_0__23_), .D(_4548__bF_buf40), .Y(_4593_) );
OAI21X1 OAI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_4592_), .B(_4547__bF_buf40), .C(_4593_), .Y(_3672__23_) );
INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__24_), .Y(_4594_) );
AOI22X1 AOI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[504]), .C(w_mem_inst_w_mem_0__24_), .D(_4548__bF_buf39), .Y(_4595_) );
OAI21X1 OAI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_4594_), .B(_4547__bF_buf39), .C(_4595_), .Y(_3672__24_) );
INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__25_), .Y(_4596_) );
AOI22X1 AOI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[505]), .C(w_mem_inst_w_mem_0__25_), .D(_4548__bF_buf38), .Y(_4597_) );
OAI21X1 OAI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_4596_), .B(_4547__bF_buf38), .C(_4597_), .Y(_3672__25_) );
INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__26_), .Y(_4598_) );
AOI22X1 AOI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[506]), .C(w_mem_inst_w_mem_0__26_), .D(_4548__bF_buf37), .Y(_4599_) );
OAI21X1 OAI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_4598_), .B(_4547__bF_buf37), .C(_4599_), .Y(_3672__26_) );
INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__27_), .Y(_4600_) );
AOI22X1 AOI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[507]), .C(w_mem_inst_w_mem_0__27_), .D(_4548__bF_buf36), .Y(_4601_) );
OAI21X1 OAI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_4600_), .B(_4547__bF_buf36), .C(_4601_), .Y(_3672__27_) );
INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__28_), .Y(_4602_) );
AOI22X1 AOI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[508]), .C(w_mem_inst_w_mem_0__28_), .D(_4548__bF_buf35), .Y(_4603_) );
OAI21X1 OAI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_4602_), .B(_4547__bF_buf35), .C(_4603_), .Y(_3672__28_) );
INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__29_), .Y(_4604_) );
AOI22X1 AOI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[509]), .C(w_mem_inst_w_mem_0__29_), .D(_4548__bF_buf34), .Y(_4605_) );
OAI21X1 OAI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_4604_), .B(_4547__bF_buf34), .C(_4605_), .Y(_3672__29_) );
INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__30_), .Y(_4606_) );
AOI22X1 AOI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[510]), .C(w_mem_inst_w_mem_0__30_), .D(_4548__bF_buf33), .Y(_4607_) );
OAI21X1 OAI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_4606_), .B(_4547__bF_buf33), .C(_4607_), .Y(_3672__30_) );
INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__31_), .Y(_4608_) );
AOI22X1 AOI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[511]), .C(w_mem_inst_w_mem_0__31_), .D(_4548__bF_buf32), .Y(_4609_) );
OAI21X1 OAI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_4608_), .B(_4547__bF_buf32), .C(_4609_), .Y(_3672__31_) );
AOI22X1 AOI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[448]), .C(w_mem_inst_w_mem_1__0_), .D(_4548__bF_buf31), .Y(_4610_) );
OAI21X1 OAI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_4547__bF_buf31), .C(_4610_), .Y(_3679__0_) );
INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__1_), .Y(_4611_) );
AOI22X1 AOI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[449]), .C(w_mem_inst_w_mem_1__1_), .D(_4548__bF_buf30), .Y(_4612_) );
OAI21X1 OAI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_4611_), .B(_4547__bF_buf30), .C(_4612_), .Y(_3679__1_) );
INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__2_), .Y(_4613_) );
AOI22X1 AOI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[450]), .C(w_mem_inst_w_mem_1__2_), .D(_4548__bF_buf29), .Y(_4614_) );
OAI21X1 OAI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_4613_), .B(_4547__bF_buf29), .C(_4614_), .Y(_3679__2_) );
INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__3_), .Y(_4615_) );
AOI22X1 AOI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[451]), .C(w_mem_inst_w_mem_1__3_), .D(_4548__bF_buf28), .Y(_4616_) );
OAI21X1 OAI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_4615_), .B(_4547__bF_buf28), .C(_4616_), .Y(_3679__3_) );
INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__4_), .Y(_4617_) );
AOI22X1 AOI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[452]), .C(w_mem_inst_w_mem_1__4_), .D(_4548__bF_buf27), .Y(_4618_) );
OAI21X1 OAI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_4617_), .B(_4547__bF_buf27), .C(_4618_), .Y(_3679__4_) );
INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__5_), .Y(_4619_) );
AOI22X1 AOI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[453]), .C(w_mem_inst_w_mem_1__5_), .D(_4548__bF_buf26), .Y(_4620_) );
OAI21X1 OAI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_4619_), .B(_4547__bF_buf26), .C(_4620_), .Y(_3679__5_) );
INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__6_), .Y(_4621_) );
AOI22X1 AOI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[454]), .C(w_mem_inst_w_mem_1__6_), .D(_4548__bF_buf25), .Y(_4622_) );
OAI21X1 OAI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_4621_), .B(_4547__bF_buf25), .C(_4622_), .Y(_3679__6_) );
INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__7_), .Y(_4623_) );
AOI22X1 AOI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[455]), .C(w_mem_inst_w_mem_1__7_), .D(_4548__bF_buf24), .Y(_4624_) );
OAI21X1 OAI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_4623_), .B(_4547__bF_buf24), .C(_4624_), .Y(_3679__7_) );
INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__8_), .Y(_4625_) );
AOI22X1 AOI22X1_136 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[456]), .C(w_mem_inst_w_mem_1__8_), .D(_4548__bF_buf23), .Y(_4626_) );
OAI21X1 OAI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_4625_), .B(_4547__bF_buf23), .C(_4626_), .Y(_3679__8_) );
AOI22X1 AOI22X1_137 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[457]), .C(w_mem_inst_w_mem_1__9_), .D(_4548__bF_buf22), .Y(_4627_) );
OAI21X1 OAI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_3960_), .B(_4547__bF_buf22), .C(_4627_), .Y(_3679__9_) );
AOI22X1 AOI22X1_138 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[458]), .C(w_mem_inst_w_mem_1__10_), .D(_4548__bF_buf21), .Y(_4628_) );
OAI21X1 OAI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3983_), .B(_4547__bF_buf21), .C(_4628_), .Y(_3679__10_) );
INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__11_), .Y(_4629_) );
AOI22X1 AOI22X1_139 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[459]), .C(w_mem_inst_w_mem_1__11_), .D(_4548__bF_buf20), .Y(_4630_) );
OAI21X1 OAI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_4629_), .B(_4547__bF_buf20), .C(_4630_), .Y(_3679__11_) );
INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__12_), .Y(_4631_) );
AOI22X1 AOI22X1_140 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[460]), .C(w_mem_inst_w_mem_1__12_), .D(_4548__bF_buf19), .Y(_4632_) );
OAI21X1 OAI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_4631_), .B(_4547__bF_buf19), .C(_4632_), .Y(_3679__12_) );
AOI22X1 AOI22X1_141 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[461]), .C(w_mem_inst_w_mem_1__13_), .D(_4548__bF_buf18), .Y(_4633_) );
OAI21X1 OAI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_4058_), .B(_4547__bF_buf18), .C(_4633_), .Y(_3679__13_) );
INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__14_), .Y(_4634_) );
AOI22X1 AOI22X1_142 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[462]), .C(w_mem_inst_w_mem_1__14_), .D(_4548__bF_buf17), .Y(_4635_) );
OAI21X1 OAI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_4634_), .B(_4547__bF_buf17), .C(_4635_), .Y(_3679__14_) );
INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__15_), .Y(_4636_) );
AOI22X1 AOI22X1_143 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[463]), .C(w_mem_inst_w_mem_1__15_), .D(_4548__bF_buf16), .Y(_4637_) );
OAI21X1 OAI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_4636_), .B(_4547__bF_buf16), .C(_4637_), .Y(_3679__15_) );
INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__16_), .Y(_4638_) );
AOI22X1 AOI22X1_144 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[464]), .C(w_mem_inst_w_mem_1__16_), .D(_4548__bF_buf15), .Y(_4639_) );
OAI21X1 OAI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_4638_), .B(_4547__bF_buf15), .C(_4639_), .Y(_3679__16_) );
AOI22X1 AOI22X1_145 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[465]), .C(w_mem_inst_w_mem_1__17_), .D(_4548__bF_buf14), .Y(_4640_) );
OAI21X1 OAI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_4158_), .B(_4547__bF_buf14), .C(_4640_), .Y(_3679__17_) );
AOI22X1 AOI22X1_146 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[466]), .C(w_mem_inst_w_mem_1__18_), .D(_4548__bF_buf13), .Y(_4641_) );
OAI21X1 OAI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_4181_), .B(_4547__bF_buf13), .C(_4641_), .Y(_3679__18_) );
INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__19_), .Y(_4642_) );
AOI22X1 AOI22X1_147 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[467]), .C(w_mem_inst_w_mem_1__19_), .D(_4548__bF_buf12), .Y(_4643_) );
OAI21X1 OAI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_4642_), .B(_4547__bF_buf12), .C(_4643_), .Y(_3679__19_) );
INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__20_), .Y(_4644_) );
AOI22X1 AOI22X1_148 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[468]), .C(w_mem_inst_w_mem_1__20_), .D(_4548__bF_buf11), .Y(_4645_) );
OAI21X1 OAI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_4644_), .B(_4547__bF_buf11), .C(_4645_), .Y(_3679__20_) );
AOI22X1 AOI22X1_149 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[469]), .C(w_mem_inst_w_mem_1__21_), .D(_4548__bF_buf10), .Y(_4646_) );
OAI21X1 OAI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_4256_), .B(_4547__bF_buf10), .C(_4646_), .Y(_3679__21_) );
INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__22_), .Y(_4647_) );
AOI22X1 AOI22X1_150 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[470]), .C(w_mem_inst_w_mem_1__22_), .D(_4548__bF_buf9), .Y(_4648_) );
OAI21X1 OAI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_4647_), .B(_4547__bF_buf9), .C(_4648_), .Y(_3679__22_) );
INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__23_), .Y(_4649_) );
AOI22X1 AOI22X1_151 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[471]), .C(w_mem_inst_w_mem_1__23_), .D(_4548__bF_buf8), .Y(_4650_) );
OAI21X1 OAI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_4649_), .B(_4547__bF_buf8), .C(_4650_), .Y(_3679__23_) );
INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__24_), .Y(_4651_) );
AOI22X1 AOI22X1_152 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[472]), .C(w_mem_inst_w_mem_1__24_), .D(_4548__bF_buf7), .Y(_4652_) );
OAI21X1 OAI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_4651_), .B(_4547__bF_buf7), .C(_4652_), .Y(_3679__24_) );
AOI22X1 AOI22X1_153 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[473]), .C(w_mem_inst_w_mem_1__25_), .D(_4548__bF_buf6), .Y(_4653_) );
OAI21X1 OAI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_4356_), .B(_4547__bF_buf6), .C(_4653_), .Y(_3679__25_) );
AOI22X1 AOI22X1_154 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[474]), .C(w_mem_inst_w_mem_1__26_), .D(_4548__bF_buf5), .Y(_4654_) );
OAI21X1 OAI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_4379_), .B(_4547__bF_buf5), .C(_4654_), .Y(_3679__26_) );
INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__27_), .Y(_4655_) );
AOI22X1 AOI22X1_155 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[475]), .C(w_mem_inst_w_mem_1__27_), .D(_4548__bF_buf4), .Y(_4656_) );
OAI21X1 OAI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_4655_), .B(_4547__bF_buf4), .C(_4656_), .Y(_3679__27_) );
INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__28_), .Y(_4657_) );
AOI22X1 AOI22X1_156 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[476]), .C(w_mem_inst_w_mem_1__28_), .D(_4548__bF_buf3), .Y(_4658_) );
OAI21X1 OAI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_4657_), .B(_4547__bF_buf3), .C(_4658_), .Y(_3679__28_) );
AOI22X1 AOI22X1_157 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[477]), .C(w_mem_inst_w_mem_1__29_), .D(_4548__bF_buf2), .Y(_4659_) );
OAI21X1 OAI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_4454_), .B(_4547__bF_buf2), .C(_4659_), .Y(_3679__29_) );
INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__30_), .Y(_4660_) );
AOI22X1 AOI22X1_158 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[478]), .C(w_mem_inst_w_mem_1__30_), .D(_4548__bF_buf1), .Y(_4661_) );
OAI21X1 OAI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_4660_), .B(_4547__bF_buf1), .C(_4661_), .Y(_3679__30_) );
INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__31_), .Y(_4662_) );
AOI22X1 AOI22X1_159 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[479]), .C(w_mem_inst_w_mem_1__31_), .D(_4548__bF_buf0), .Y(_4663_) );
OAI21X1 OAI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_4662_), .B(_4547__bF_buf0), .C(_4663_), .Y(_3679__31_) );
INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__0_), .Y(_4664_) );
AOI22X1 AOI22X1_160 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[416]), .C(w_mem_inst_w_mem_2__0_), .D(_4548__bF_buf63), .Y(_4665_) );
OAI21X1 OAI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_4664_), .B(_4547__bF_buf63), .C(_4665_), .Y(_3680__0_) );
AOI22X1 AOI22X1_161 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[417]), .C(w_mem_inst_w_mem_2__1_), .D(_4548__bF_buf62), .Y(_4666_) );
OAI21X1 OAI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_3762_), .B(_4547__bF_buf62), .C(_4666_), .Y(_3680__1_) );
INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__2_), .Y(_4667_) );
AOI22X1 AOI22X1_162 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[418]), .C(w_mem_inst_w_mem_2__2_), .D(_4548__bF_buf61), .Y(_4668_) );
OAI21X1 OAI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_4667_), .B(_4547__bF_buf61), .C(_4668_), .Y(_3680__2_) );
AOI22X1 AOI22X1_163 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[419]), .C(w_mem_inst_w_mem_2__3_), .D(_4548__bF_buf60), .Y(_4669_) );
OAI21X1 OAI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3814_), .B(_4547__bF_buf60), .C(_4669_), .Y(_3680__3_) );
INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__4_), .Y(_4670_) );
AOI22X1 AOI22X1_164 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[420]), .C(w_mem_inst_w_mem_2__4_), .D(_4548__bF_buf59), .Y(_4671_) );
OAI21X1 OAI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_4670_), .B(_4547__bF_buf59), .C(_4671_), .Y(_3680__4_) );
INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__5_), .Y(_4672_) );
AOI22X1 AOI22X1_165 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[421]), .C(w_mem_inst_w_mem_2__5_), .D(_4548__bF_buf58), .Y(_4673_) );
OAI21X1 OAI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_4672_), .B(_4547__bF_buf58), .C(_4673_), .Y(_3680__5_) );
INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__6_), .Y(_4674_) );
AOI22X1 AOI22X1_166 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[422]), .C(w_mem_inst_w_mem_2__6_), .D(_4548__bF_buf57), .Y(_4675_) );
OAI21X1 OAI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_4674_), .B(_4547__bF_buf57), .C(_4675_), .Y(_3680__6_) );
INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__7_), .Y(_4676_) );
AOI22X1 AOI22X1_167 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[423]), .C(w_mem_inst_w_mem_2__7_), .D(_4548__bF_buf56), .Y(_4677_) );
OAI21X1 OAI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_4676_), .B(_4547__bF_buf56), .C(_4677_), .Y(_3680__7_) );
AOI22X1 AOI22X1_168 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[424]), .C(w_mem_inst_w_mem_2__8_), .D(_4548__bF_buf55), .Y(_4678_) );
OAI21X1 OAI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_3939_), .B(_4547__bF_buf55), .C(_4678_), .Y(_3680__8_) );
AOI22X1 AOI22X1_169 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[425]), .C(w_mem_inst_w_mem_2__9_), .D(_4548__bF_buf54), .Y(_4679_) );
OAI21X1 OAI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_3958_), .B(_4547__bF_buf54), .C(_4679_), .Y(_3680__9_) );
INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__10_), .Y(_4680_) );
AOI22X1 AOI22X1_170 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[426]), .C(w_mem_inst_w_mem_2__10_), .D(_4548__bF_buf53), .Y(_4681_) );
OAI21X1 OAI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_4680_), .B(_4547__bF_buf53), .C(_4681_), .Y(_3680__10_) );
INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__11_), .Y(_4682_) );
AOI22X1 AOI22X1_171 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[427]), .C(w_mem_inst_w_mem_2__11_), .D(_4548__bF_buf52), .Y(_4683_) );
OAI21X1 OAI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_4682_), .B(_4547__bF_buf52), .C(_4683_), .Y(_3680__11_) );
INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__12_), .Y(_4684_) );
AOI22X1 AOI22X1_172 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[428]), .C(w_mem_inst_w_mem_2__12_), .D(_4548__bF_buf51), .Y(_4685_) );
OAI21X1 OAI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_4684_), .B(_4547__bF_buf51), .C(_4685_), .Y(_3680__12_) );
INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__13_), .Y(_4686_) );
AOI22X1 AOI22X1_173 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[429]), .C(w_mem_inst_w_mem_2__13_), .D(_4548__bF_buf50), .Y(_4687_) );
OAI21X1 OAI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_4686_), .B(_4547__bF_buf50), .C(_4687_), .Y(_3680__13_) );
INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__14_), .Y(_4688_) );
AOI22X1 AOI22X1_174 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[430]), .C(w_mem_inst_w_mem_2__14_), .D(_4548__bF_buf49), .Y(_4689_) );
OAI21X1 OAI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_4688_), .B(_4547__bF_buf49), .C(_4689_), .Y(_3680__14_) );
INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__15_), .Y(_4690_) );
AOI22X1 AOI22X1_175 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[431]), .C(w_mem_inst_w_mem_2__15_), .D(_4548__bF_buf48), .Y(_4691_) );
OAI21X1 OAI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_4690_), .B(_4547__bF_buf48), .C(_4691_), .Y(_3680__15_) );
AOI22X1 AOI22X1_176 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[432]), .C(w_mem_inst_w_mem_2__16_), .D(_4548__bF_buf47), .Y(_4692_) );
OAI21X1 OAI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_4137_), .B(_4547__bF_buf47), .C(_4692_), .Y(_3680__16_) );
AOI22X1 AOI22X1_177 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[433]), .C(w_mem_inst_w_mem_2__17_), .D(_4548__bF_buf46), .Y(_4693_) );
OAI21X1 OAI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_4156_), .B(_4547__bF_buf46), .C(_4693_), .Y(_3680__17_) );
INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__18_), .Y(_4694_) );
AOI22X1 AOI22X1_178 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[434]), .C(w_mem_inst_w_mem_2__18_), .D(_4548__bF_buf45), .Y(_4695_) );
OAI21X1 OAI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_4694_), .B(_4547__bF_buf45), .C(_4695_), .Y(_3680__18_) );
INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__19_), .Y(_4696_) );
AOI22X1 AOI22X1_179 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[435]), .C(w_mem_inst_w_mem_2__19_), .D(_4548__bF_buf44), .Y(_4697_) );
OAI21X1 OAI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_4696_), .B(_4547__bF_buf44), .C(_4697_), .Y(_3680__19_) );
INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__20_), .Y(_4698_) );
AOI22X1 AOI22X1_180 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[436]), .C(w_mem_inst_w_mem_2__20_), .D(_4548__bF_buf43), .Y(_4699_) );
OAI21X1 OAI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_4698_), .B(_4547__bF_buf43), .C(_4699_), .Y(_3680__20_) );
INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__21_), .Y(_4700_) );
AOI22X1 AOI22X1_181 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[437]), .C(w_mem_inst_w_mem_2__21_), .D(_4548__bF_buf42), .Y(_4701_) );
OAI21X1 OAI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_4700_), .B(_4547__bF_buf42), .C(_4701_), .Y(_3680__21_) );
INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__22_), .Y(_4702_) );
AOI22X1 AOI22X1_182 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[438]), .C(w_mem_inst_w_mem_2__22_), .D(_4548__bF_buf41), .Y(_4703_) );
OAI21X1 OAI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_4702_), .B(_4547__bF_buf41), .C(_4703_), .Y(_3680__22_) );
INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__23_), .Y(_4704_) );
AOI22X1 AOI22X1_183 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[439]), .C(w_mem_inst_w_mem_2__23_), .D(_4548__bF_buf40), .Y(_4705_) );
OAI21X1 OAI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_4704_), .B(_4547__bF_buf40), .C(_4705_), .Y(_3680__23_) );
AOI22X1 AOI22X1_184 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[440]), .C(w_mem_inst_w_mem_2__24_), .D(_4548__bF_buf39), .Y(_4706_) );
OAI21X1 OAI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_4335_), .B(_4547__bF_buf39), .C(_4706_), .Y(_3680__24_) );
AOI22X1 AOI22X1_185 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[441]), .C(w_mem_inst_w_mem_2__25_), .D(_4548__bF_buf38), .Y(_4707_) );
OAI21X1 OAI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_4354_), .B(_4547__bF_buf38), .C(_4707_), .Y(_3680__25_) );
INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__26_), .Y(_4708_) );
AOI22X1 AOI22X1_186 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[442]), .C(w_mem_inst_w_mem_2__26_), .D(_4548__bF_buf37), .Y(_4709_) );
OAI21X1 OAI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_4708_), .B(_4547__bF_buf37), .C(_4709_), .Y(_3680__26_) );
INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__27_), .Y(_4710_) );
AOI22X1 AOI22X1_187 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[443]), .C(w_mem_inst_w_mem_2__27_), .D(_4548__bF_buf36), .Y(_4711_) );
OAI21X1 OAI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_4710_), .B(_4547__bF_buf36), .C(_4711_), .Y(_3680__27_) );
INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__28_), .Y(_4712_) );
AOI22X1 AOI22X1_188 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[444]), .C(w_mem_inst_w_mem_2__28_), .D(_4548__bF_buf35), .Y(_4713_) );
OAI21X1 OAI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_4712_), .B(_4547__bF_buf35), .C(_4713_), .Y(_3680__28_) );
INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__29_), .Y(_4714_) );
AOI22X1 AOI22X1_189 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[445]), .C(w_mem_inst_w_mem_2__29_), .D(_4548__bF_buf34), .Y(_4715_) );
OAI21X1 OAI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_4714_), .B(_4547__bF_buf34), .C(_4715_), .Y(_3680__29_) );
INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__30_), .Y(_4716_) );
AOI22X1 AOI22X1_190 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[446]), .C(w_mem_inst_w_mem_2__30_), .D(_4548__bF_buf33), .Y(_4717_) );
OAI21X1 OAI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_4716_), .B(_4547__bF_buf33), .C(_4717_), .Y(_3680__30_) );
INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__31_), .Y(_4718_) );
AOI22X1 AOI22X1_191 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[447]), .C(w_mem_inst_w_mem_2__31_), .D(_4548__bF_buf32), .Y(_4719_) );
OAI21X1 OAI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_4718_), .B(_4547__bF_buf32), .C(_4719_), .Y(_3680__31_) );
INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__0_), .Y(_4720_) );
AOI22X1 AOI22X1_192 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[384]), .C(w_mem_inst_w_mem_3__0_), .D(_4548__bF_buf31), .Y(_4721_) );
OAI21X1 OAI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_4720_), .B(_4547__bF_buf31), .C(_4721_), .Y(_3681__0_) );
INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__1_), .Y(_4722_) );
AOI22X1 AOI22X1_193 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[385]), .C(w_mem_inst_w_mem_3__1_), .D(_4548__bF_buf30), .Y(_4723_) );
OAI21X1 OAI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_4722_), .B(_4547__bF_buf30), .C(_4723_), .Y(_3681__1_) );
INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__2_), .Y(_4724_) );
AOI22X1 AOI22X1_194 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[386]), .C(w_mem_inst_w_mem_3__2_), .D(_4548__bF_buf29), .Y(_4725_) );
OAI21X1 OAI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_4724_), .B(_4547__bF_buf29), .C(_4725_), .Y(_3681__2_) );
INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__3_), .Y(_4726_) );
AOI22X1 AOI22X1_195 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[387]), .C(w_mem_inst_w_mem_3__3_), .D(_4548__bF_buf28), .Y(_4727_) );
OAI21X1 OAI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_4726_), .B(_4547__bF_buf28), .C(_4727_), .Y(_3681__3_) );
AOI22X1 AOI22X1_196 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[388]), .C(w_mem_inst_w_mem_3__4_), .D(_4548__bF_buf27), .Y(_4728_) );
OAI21X1 OAI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_3832_), .B(_4547__bF_buf27), .C(_4728_), .Y(_3681__4_) );
INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__5_), .Y(_4729_) );
AOI22X1 AOI22X1_197 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[389]), .C(w_mem_inst_w_mem_3__5_), .D(_4548__bF_buf26), .Y(_4730_) );
OAI21X1 OAI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_4729_), .B(_4547__bF_buf26), .C(_4730_), .Y(_3681__5_) );
INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__6_), .Y(_4731_) );
AOI22X1 AOI22X1_198 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[390]), .C(w_mem_inst_w_mem_3__6_), .D(_4548__bF_buf25), .Y(_4732_) );
OAI21X1 OAI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_4731_), .B(_4547__bF_buf25), .C(_4732_), .Y(_3681__6_) );
AOI22X1 AOI22X1_199 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[391]), .C(w_mem_inst_w_mem_3__7_), .D(_4548__bF_buf24), .Y(_4733_) );
OAI21X1 OAI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_3909_), .B(_4547__bF_buf24), .C(_4733_), .Y(_3681__7_) );
INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__8_), .Y(_4734_) );
AOI22X1 AOI22X1_200 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[392]), .C(w_mem_inst_w_mem_3__8_), .D(_4548__bF_buf23), .Y(_4735_) );
OAI21X1 OAI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_4734_), .B(_4547__bF_buf23), .C(_4735_), .Y(_3681__8_) );
INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__9_), .Y(_4736_) );
AOI22X1 AOI22X1_201 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[393]), .C(w_mem_inst_w_mem_3__9_), .D(_4548__bF_buf22), .Y(_4737_) );
OAI21X1 OAI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_4736_), .B(_4547__bF_buf22), .C(_4737_), .Y(_3681__9_) );
INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__10_), .Y(_4738_) );
AOI22X1 AOI22X1_202 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[394]), .C(w_mem_inst_w_mem_3__10_), .D(_4548__bF_buf21), .Y(_4739_) );
OAI21X1 OAI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_4738_), .B(_4547__bF_buf21), .C(_4739_), .Y(_3681__10_) );
AOI22X1 AOI22X1_203 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[395]), .C(w_mem_inst_w_mem_3__11_), .D(_4548__bF_buf20), .Y(_4740_) );
OAI21X1 OAI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_4008_), .B(_4547__bF_buf20), .C(_4740_), .Y(_3681__11_) );
AOI22X1 AOI22X1_204 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[396]), .C(w_mem_inst_w_mem_3__12_), .D(_4548__bF_buf19), .Y(_4741_) );
OAI21X1 OAI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_4033_), .B(_4547__bF_buf19), .C(_4741_), .Y(_3681__12_) );
INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__13_), .Y(_4742_) );
AOI22X1 AOI22X1_205 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[397]), .C(w_mem_inst_w_mem_3__13_), .D(_4548__bF_buf18), .Y(_4743_) );
OAI21X1 OAI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_4742_), .B(_4547__bF_buf18), .C(_4743_), .Y(_3681__13_) );
INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__14_), .Y(_4744_) );
AOI22X1 AOI22X1_206 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[398]), .C(w_mem_inst_w_mem_3__14_), .D(_4548__bF_buf17), .Y(_4745_) );
OAI21X1 OAI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_4744_), .B(_4547__bF_buf17), .C(_4745_), .Y(_3681__14_) );
AOI22X1 AOI22X1_207 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[399]), .C(w_mem_inst_w_mem_3__15_), .D(_4548__bF_buf16), .Y(_4746_) );
OAI21X1 OAI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_4107_), .B(_4547__bF_buf16), .C(_4746_), .Y(_3681__15_) );
INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__16_), .Y(_4747_) );
AOI22X1 AOI22X1_208 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[400]), .C(w_mem_inst_w_mem_3__16_), .D(_4548__bF_buf15), .Y(_4748_) );
OAI21X1 OAI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_4747_), .B(_4547__bF_buf15), .C(_4748_), .Y(_3681__16_) );
INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__17_), .Y(_4749_) );
AOI22X1 AOI22X1_209 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[401]), .C(w_mem_inst_w_mem_3__17_), .D(_4548__bF_buf14), .Y(_4750_) );
OAI21X1 OAI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_4749_), .B(_4547__bF_buf14), .C(_4750_), .Y(_3681__17_) );
INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__18_), .Y(_4751_) );
AOI22X1 AOI22X1_210 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[402]), .C(w_mem_inst_w_mem_3__18_), .D(_4548__bF_buf13), .Y(_4752_) );
OAI21X1 OAI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_4751_), .B(_4547__bF_buf13), .C(_4752_), .Y(_3681__18_) );
AOI22X1 AOI22X1_211 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[403]), .C(w_mem_inst_w_mem_3__19_), .D(_4548__bF_buf12), .Y(_4753_) );
OAI21X1 OAI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_4206_), .B(_4547__bF_buf12), .C(_4753_), .Y(_3681__19_) );
AOI22X1 AOI22X1_212 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[404]), .C(w_mem_inst_w_mem_3__20_), .D(_4548__bF_buf11), .Y(_4754_) );
OAI21X1 OAI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_4231_), .B(_4547__bF_buf11), .C(_4754_), .Y(_3681__20_) );
INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__21_), .Y(_4755_) );
AOI22X1 AOI22X1_213 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[405]), .C(w_mem_inst_w_mem_3__21_), .D(_4548__bF_buf10), .Y(_4756_) );
OAI21X1 OAI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_4755_), .B(_4547__bF_buf10), .C(_4756_), .Y(_3681__21_) );
INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__22_), .Y(_4757_) );
AOI22X1 AOI22X1_214 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[406]), .C(w_mem_inst_w_mem_3__22_), .D(_4548__bF_buf9), .Y(_4758_) );
OAI21X1 OAI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_4757_), .B(_4547__bF_buf9), .C(_4758_), .Y(_3681__22_) );
AOI22X1 AOI22X1_215 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[407]), .C(w_mem_inst_w_mem_3__23_), .D(_4548__bF_buf8), .Y(_4759_) );
OAI21X1 OAI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_4305_), .B(_4547__bF_buf8), .C(_4759_), .Y(_3681__23_) );
INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__24_), .Y(_4760_) );
AOI22X1 AOI22X1_216 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[408]), .C(w_mem_inst_w_mem_3__24_), .D(_4548__bF_buf7), .Y(_4761_) );
OAI21X1 OAI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_4760_), .B(_4547__bF_buf7), .C(_4761_), .Y(_3681__24_) );
INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__25_), .Y(_4762_) );
AOI22X1 AOI22X1_217 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[409]), .C(w_mem_inst_w_mem_3__25_), .D(_4548__bF_buf6), .Y(_4763_) );
OAI21X1 OAI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_4762_), .B(_4547__bF_buf6), .C(_4763_), .Y(_3681__25_) );
INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__26_), .Y(_4764_) );
AOI22X1 AOI22X1_218 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[410]), .C(w_mem_inst_w_mem_3__26_), .D(_4548__bF_buf5), .Y(_4765_) );
OAI21X1 OAI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_4764_), .B(_4547__bF_buf5), .C(_4765_), .Y(_3681__26_) );
AOI22X1 AOI22X1_219 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[411]), .C(w_mem_inst_w_mem_3__27_), .D(_4548__bF_buf4), .Y(_4766_) );
OAI21X1 OAI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_4404_), .B(_4547__bF_buf4), .C(_4766_), .Y(_3681__27_) );
AOI22X1 AOI22X1_220 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[412]), .C(w_mem_inst_w_mem_3__28_), .D(_4548__bF_buf3), .Y(_4767_) );
OAI21X1 OAI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_4429_), .B(_4547__bF_buf3), .C(_4767_), .Y(_3681__28_) );
INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__29_), .Y(_4768_) );
AOI22X1 AOI22X1_221 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[413]), .C(w_mem_inst_w_mem_3__29_), .D(_4548__bF_buf2), .Y(_4769_) );
OAI21X1 OAI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_4768_), .B(_4547__bF_buf2), .C(_4769_), .Y(_3681__29_) );
INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__30_), .Y(_4770_) );
AOI22X1 AOI22X1_222 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[414]), .C(w_mem_inst_w_mem_3__30_), .D(_4548__bF_buf1), .Y(_4771_) );
OAI21X1 OAI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_4770_), .B(_4547__bF_buf1), .C(_4771_), .Y(_3681__30_) );
AOI22X1 AOI22X1_223 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[415]), .C(w_mem_inst_w_mem_3__31_), .D(_4548__bF_buf0), .Y(_4772_) );
OAI21X1 OAI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_4503_), .B(_4547__bF_buf0), .C(_4772_), .Y(_3681__31_) );
INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__0_), .Y(_4773_) );
AOI22X1 AOI22X1_224 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[352]), .C(w_mem_inst_w_mem_4__0_), .D(_4548__bF_buf63), .Y(_4774_) );
OAI21X1 OAI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_4773_), .B(_4547__bF_buf63), .C(_4774_), .Y(_3682__0_) );
AOI22X1 AOI22X1_225 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[353]), .C(w_mem_inst_w_mem_4__1_), .D(_4548__bF_buf62), .Y(_4775_) );
OAI21X1 OAI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_4547__bF_buf62), .C(_4775_), .Y(_3682__1_) );
AOI22X1 AOI22X1_226 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[354]), .C(w_mem_inst_w_mem_4__2_), .D(_4548__bF_buf61), .Y(_4776_) );
OAI21X1 OAI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_3793_), .B(_4547__bF_buf61), .C(_4776_), .Y(_3682__2_) );
INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__3_), .Y(_4777_) );
AOI22X1 AOI22X1_227 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[355]), .C(w_mem_inst_w_mem_4__3_), .D(_4548__bF_buf60), .Y(_4778_) );
OAI21X1 OAI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_4777_), .B(_4547__bF_buf60), .C(_4778_), .Y(_3682__3_) );
AOI22X1 AOI22X1_228 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[356]), .C(w_mem_inst_w_mem_4__4_), .D(_4548__bF_buf59), .Y(_4779_) );
OAI21X1 OAI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_3841_), .B(_4547__bF_buf59), .C(_4779_), .Y(_3682__4_) );
INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__5_), .Y(_4780_) );
AOI22X1 AOI22X1_229 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[357]), .C(w_mem_inst_w_mem_4__5_), .D(_4548__bF_buf58), .Y(_4781_) );
OAI21X1 OAI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_4780_), .B(_4547__bF_buf58), .C(_4781_), .Y(_3682__5_) );
AOI22X1 AOI22X1_230 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[358]), .C(w_mem_inst_w_mem_4__6_), .D(_4548__bF_buf57), .Y(_4782_) );
OAI21X1 OAI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_3891_), .B(_4547__bF_buf57), .C(_4782_), .Y(_3682__6_) );
INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__7_), .Y(_4783_) );
AOI22X1 AOI22X1_231 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[359]), .C(w_mem_inst_w_mem_4__7_), .D(_4548__bF_buf56), .Y(_4784_) );
OAI21X1 OAI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_4783_), .B(_4547__bF_buf56), .C(_4784_), .Y(_3682__7_) );
INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__8_), .Y(_4785_) );
AOI22X1 AOI22X1_232 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[360]), .C(w_mem_inst_w_mem_4__8_), .D(_4548__bF_buf55), .Y(_4786_) );
OAI21X1 OAI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_4785_), .B(_4547__bF_buf55), .C(_4786_), .Y(_3682__8_) );
AOI22X1 AOI22X1_233 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[361]), .C(w_mem_inst_w_mem_4__9_), .D(_4548__bF_buf54), .Y(_4787_) );
OAI21X1 OAI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_3961_), .B(_4547__bF_buf54), .C(_4787_), .Y(_3682__9_) );
AOI22X1 AOI22X1_234 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[362]), .C(w_mem_inst_w_mem_4__10_), .D(_4548__bF_buf53), .Y(_4788_) );
OAI21X1 OAI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_3985_), .B(_4547__bF_buf53), .C(_4788_), .Y(_3682__10_) );
INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__11_), .Y(_4789_) );
AOI22X1 AOI22X1_235 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[363]), .C(w_mem_inst_w_mem_4__11_), .D(_4548__bF_buf52), .Y(_4790_) );
OAI21X1 OAI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_4789_), .B(_4547__bF_buf52), .C(_4790_), .Y(_3682__11_) );
AOI22X1 AOI22X1_236 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[364]), .C(w_mem_inst_w_mem_4__12_), .D(_4548__bF_buf51), .Y(_4791_) );
OAI21X1 OAI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_4039_), .B(_4547__bF_buf51), .C(_4791_), .Y(_3682__12_) );
INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__13_), .Y(_4792_) );
AOI22X1 AOI22X1_237 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[365]), .C(w_mem_inst_w_mem_4__13_), .D(_4548__bF_buf50), .Y(_4793_) );
OAI21X1 OAI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_4792_), .B(_4547__bF_buf50), .C(_4793_), .Y(_3682__13_) );
AOI22X1 AOI22X1_238 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[366]), .C(w_mem_inst_w_mem_4__14_), .D(_4548__bF_buf49), .Y(_4794_) );
OAI21X1 OAI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_4089_), .B(_4547__bF_buf49), .C(_4794_), .Y(_3682__14_) );
INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__15_), .Y(_4795_) );
AOI22X1 AOI22X1_239 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[367]), .C(w_mem_inst_w_mem_4__15_), .D(_4548__bF_buf48), .Y(_4796_) );
OAI21X1 OAI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_4795_), .B(_4547__bF_buf48), .C(_4796_), .Y(_3682__15_) );
INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__16_), .Y(_4797_) );
AOI22X1 AOI22X1_240 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[368]), .C(w_mem_inst_w_mem_4__16_), .D(_4548__bF_buf47), .Y(_4798_) );
OAI21X1 OAI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_4797_), .B(_4547__bF_buf47), .C(_4798_), .Y(_3682__16_) );
AOI22X1 AOI22X1_241 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[369]), .C(w_mem_inst_w_mem_4__17_), .D(_4548__bF_buf46), .Y(_4799_) );
OAI21X1 OAI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_4159_), .B(_4547__bF_buf46), .C(_4799_), .Y(_3682__17_) );
AOI22X1 AOI22X1_242 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[370]), .C(w_mem_inst_w_mem_4__18_), .D(_4548__bF_buf45), .Y(_4800_) );
OAI21X1 OAI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_4183_), .B(_4547__bF_buf45), .C(_4800_), .Y(_3682__18_) );
INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__19_), .Y(_4801_) );
AOI22X1 AOI22X1_243 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[371]), .C(w_mem_inst_w_mem_4__19_), .D(_4548__bF_buf44), .Y(_4802_) );
OAI21X1 OAI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_4801_), .B(_4547__bF_buf44), .C(_4802_), .Y(_3682__19_) );
AOI22X1 AOI22X1_244 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[372]), .C(w_mem_inst_w_mem_4__20_), .D(_4548__bF_buf43), .Y(_4803_) );
OAI21X1 OAI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_4237_), .B(_4547__bF_buf43), .C(_4803_), .Y(_3682__20_) );
INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__21_), .Y(_4804_) );
AOI22X1 AOI22X1_245 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[373]), .C(w_mem_inst_w_mem_4__21_), .D(_4548__bF_buf42), .Y(_4805_) );
OAI21X1 OAI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_4804_), .B(_4547__bF_buf42), .C(_4805_), .Y(_3682__21_) );
AOI22X1 AOI22X1_246 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[374]), .C(w_mem_inst_w_mem_4__22_), .D(_4548__bF_buf41), .Y(_4806_) );
OAI21X1 OAI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_4287_), .B(_4547__bF_buf41), .C(_4806_), .Y(_3682__22_) );
INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__23_), .Y(_4807_) );
AOI22X1 AOI22X1_247 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[375]), .C(w_mem_inst_w_mem_4__23_), .D(_4548__bF_buf40), .Y(_4808_) );
OAI21X1 OAI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_4807_), .B(_4547__bF_buf40), .C(_4808_), .Y(_3682__23_) );
INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__24_), .Y(_4809_) );
AOI22X1 AOI22X1_248 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[376]), .C(w_mem_inst_w_mem_4__24_), .D(_4548__bF_buf39), .Y(_4810_) );
OAI21X1 OAI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_4809_), .B(_4547__bF_buf39), .C(_4810_), .Y(_3682__24_) );
AOI22X1 AOI22X1_249 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[377]), .C(w_mem_inst_w_mem_4__25_), .D(_4548__bF_buf38), .Y(_4811_) );
OAI21X1 OAI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_4357_), .B(_4547__bF_buf38), .C(_4811_), .Y(_3682__25_) );
AOI22X1 AOI22X1_250 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[378]), .C(w_mem_inst_w_mem_4__26_), .D(_4548__bF_buf37), .Y(_4812_) );
OAI21X1 OAI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_4381_), .B(_4547__bF_buf37), .C(_4812_), .Y(_3682__26_) );
INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__27_), .Y(_4813_) );
AOI22X1 AOI22X1_251 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[379]), .C(w_mem_inst_w_mem_4__27_), .D(_4548__bF_buf36), .Y(_4814_) );
OAI21X1 OAI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_4813_), .B(_4547__bF_buf36), .C(_4814_), .Y(_3682__27_) );
AOI22X1 AOI22X1_252 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[380]), .C(w_mem_inst_w_mem_4__28_), .D(_4548__bF_buf35), .Y(_4815_) );
OAI21X1 OAI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_4435_), .B(_4547__bF_buf35), .C(_4815_), .Y(_3682__28_) );
INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__29_), .Y(_4816_) );
AOI22X1 AOI22X1_253 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[381]), .C(w_mem_inst_w_mem_4__29_), .D(_4548__bF_buf34), .Y(_4817_) );
OAI21X1 OAI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_4816_), .B(_4547__bF_buf34), .C(_4817_), .Y(_3682__29_) );
AOI22X1 AOI22X1_254 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[382]), .C(w_mem_inst_w_mem_4__30_), .D(_4548__bF_buf33), .Y(_4818_) );
OAI21X1 OAI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_4485_), .B(_4547__bF_buf33), .C(_4818_), .Y(_3682__30_) );
INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__31_), .Y(_4819_) );
AOI22X1 AOI22X1_255 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[383]), .C(w_mem_inst_w_mem_4__31_), .D(_4548__bF_buf32), .Y(_4820_) );
OAI21X1 OAI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_4819_), .B(_4547__bF_buf32), .C(_4820_), .Y(_3682__31_) );
AOI22X1 AOI22X1_256 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[320]), .C(w_mem_inst_w_mem_5__0_), .D(_4548__bF_buf31), .Y(_4821_) );
OAI21X1 OAI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_4547__bF_buf31), .C(_4821_), .Y(_3683__0_) );
INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__1_), .Y(_4822_) );
AOI22X1 AOI22X1_257 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[321]), .C(w_mem_inst_w_mem_5__1_), .D(_4548__bF_buf30), .Y(_4823_) );
OAI21X1 OAI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_4822_), .B(_4547__bF_buf30), .C(_4823_), .Y(_3683__1_) );
INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__2_), .Y(_4824_) );
AOI22X1 AOI22X1_258 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[322]), .C(w_mem_inst_w_mem_5__2_), .D(_4548__bF_buf29), .Y(_4825_) );
OAI21X1 OAI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_4824_), .B(_4547__bF_buf29), .C(_4825_), .Y(_3683__2_) );
INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__3_), .Y(_4826_) );
AOI22X1 AOI22X1_259 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[323]), .C(w_mem_inst_w_mem_5__3_), .D(_4548__bF_buf28), .Y(_4827_) );
OAI21X1 OAI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_4826_), .B(_4547__bF_buf28), .C(_4827_), .Y(_3683__3_) );
INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__4_), .Y(_4828_) );
AOI22X1 AOI22X1_260 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[324]), .C(w_mem_inst_w_mem_5__4_), .D(_4548__bF_buf27), .Y(_4829_) );
OAI21X1 OAI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_4828_), .B(_4547__bF_buf27), .C(_4829_), .Y(_3683__4_) );
INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__5_), .Y(_4830_) );
AOI22X1 AOI22X1_261 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[325]), .C(w_mem_inst_w_mem_5__5_), .D(_4548__bF_buf26), .Y(_4831_) );
OAI21X1 OAI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_4830_), .B(_4547__bF_buf26), .C(_4831_), .Y(_3683__5_) );
INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__6_), .Y(_4832_) );
AOI22X1 AOI22X1_262 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[326]), .C(w_mem_inst_w_mem_5__6_), .D(_4548__bF_buf25), .Y(_4833_) );
OAI21X1 OAI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_4832_), .B(_4547__bF_buf25), .C(_4833_), .Y(_3683__6_) );
AOI22X1 AOI22X1_263 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[327]), .C(w_mem_inst_w_mem_5__7_), .D(_4548__bF_buf24), .Y(_4834_) );
OAI21X1 OAI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_3914_), .B(_4547__bF_buf24), .C(_4834_), .Y(_3683__7_) );
AOI22X1 AOI22X1_264 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[328]), .C(w_mem_inst_w_mem_5__8_), .D(_4548__bF_buf23), .Y(_4835_) );
OAI21X1 OAI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_3933_), .B(_4547__bF_buf23), .C(_4835_), .Y(_3683__8_) );
INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__9_), .Y(_4836_) );
AOI22X1 AOI22X1_265 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[329]), .C(w_mem_inst_w_mem_5__9_), .D(_4548__bF_buf22), .Y(_4837_) );
OAI21X1 OAI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_4836_), .B(_4547__bF_buf22), .C(_4837_), .Y(_3683__9_) );
INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__10_), .Y(_4838_) );
AOI22X1 AOI22X1_266 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[330]), .C(w_mem_inst_w_mem_5__10_), .D(_4548__bF_buf21), .Y(_4839_) );
OAI21X1 OAI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_4838_), .B(_4547__bF_buf21), .C(_4839_), .Y(_3683__10_) );
AOI22X1 AOI22X1_267 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[331]), .C(w_mem_inst_w_mem_5__11_), .D(_4548__bF_buf20), .Y(_4840_) );
OAI21X1 OAI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_4010_), .B(_4547__bF_buf20), .C(_4840_), .Y(_3683__11_) );
INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__12_), .Y(_4841_) );
AOI22X1 AOI22X1_268 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[332]), .C(w_mem_inst_w_mem_5__12_), .D(_4548__bF_buf19), .Y(_4842_) );
OAI21X1 OAI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_4841_), .B(_4547__bF_buf19), .C(_4842_), .Y(_3683__12_) );
AOI22X1 AOI22X1_269 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[333]), .C(w_mem_inst_w_mem_5__13_), .D(_4548__bF_buf18), .Y(_4843_) );
OAI21X1 OAI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_4060_), .B(_4547__bF_buf18), .C(_4843_), .Y(_3683__13_) );
INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__14_), .Y(_4844_) );
AOI22X1 AOI22X1_270 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[334]), .C(w_mem_inst_w_mem_5__14_), .D(_4548__bF_buf17), .Y(_4845_) );
OAI21X1 OAI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_4844_), .B(_4547__bF_buf17), .C(_4845_), .Y(_3683__14_) );
AOI22X1 AOI22X1_271 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[335]), .C(w_mem_inst_w_mem_5__15_), .D(_4548__bF_buf16), .Y(_4846_) );
OAI21X1 OAI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_4112_), .B(_4547__bF_buf16), .C(_4846_), .Y(_3683__15_) );
AOI22X1 AOI22X1_272 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[336]), .C(w_mem_inst_w_mem_5__16_), .D(_4548__bF_buf15), .Y(_4847_) );
OAI21X1 OAI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_4131_), .B(_4547__bF_buf15), .C(_4847_), .Y(_3683__16_) );
INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__17_), .Y(_4848_) );
AOI22X1 AOI22X1_273 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[337]), .C(w_mem_inst_w_mem_5__17_), .D(_4548__bF_buf14), .Y(_4849_) );
OAI21X1 OAI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_4848_), .B(_4547__bF_buf14), .C(_4849_), .Y(_3683__17_) );
INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__18_), .Y(_4850_) );
AOI22X1 AOI22X1_274 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[338]), .C(w_mem_inst_w_mem_5__18_), .D(_4548__bF_buf13), .Y(_4851_) );
OAI21X1 OAI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_4850_), .B(_4547__bF_buf13), .C(_4851_), .Y(_3683__18_) );
AOI22X1 AOI22X1_275 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[339]), .C(w_mem_inst_w_mem_5__19_), .D(_4548__bF_buf12), .Y(_4852_) );
OAI21X1 OAI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_4208_), .B(_4547__bF_buf12), .C(_4852_), .Y(_3683__19_) );
INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__20_), .Y(_4853_) );
AOI22X1 AOI22X1_276 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[340]), .C(w_mem_inst_w_mem_5__20_), .D(_4548__bF_buf11), .Y(_4854_) );
OAI21X1 OAI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_4853_), .B(_4547__bF_buf11), .C(_4854_), .Y(_3683__20_) );
AOI22X1 AOI22X1_277 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[341]), .C(w_mem_inst_w_mem_5__21_), .D(_4548__bF_buf10), .Y(_4855_) );
OAI21X1 OAI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_4258_), .B(_4547__bF_buf10), .C(_4855_), .Y(_3683__21_) );
INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__22_), .Y(_4856_) );
AOI22X1 AOI22X1_278 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[342]), .C(w_mem_inst_w_mem_5__22_), .D(_4548__bF_buf9), .Y(_4857_) );
OAI21X1 OAI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_4856_), .B(_4547__bF_buf9), .C(_4857_), .Y(_3683__22_) );
AOI22X1 AOI22X1_279 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[343]), .C(w_mem_inst_w_mem_5__23_), .D(_4548__bF_buf8), .Y(_4858_) );
OAI21X1 OAI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_4310_), .B(_4547__bF_buf8), .C(_4858_), .Y(_3683__23_) );
AOI22X1 AOI22X1_280 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[344]), .C(w_mem_inst_w_mem_5__24_), .D(_4548__bF_buf7), .Y(_4859_) );
OAI21X1 OAI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_4329_), .B(_4547__bF_buf7), .C(_4859_), .Y(_3683__24_) );
INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__25_), .Y(_4860_) );
AOI22X1 AOI22X1_281 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[345]), .C(w_mem_inst_w_mem_5__25_), .D(_4548__bF_buf6), .Y(_4861_) );
OAI21X1 OAI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_4860_), .B(_4547__bF_buf6), .C(_4861_), .Y(_3683__25_) );
INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__26_), .Y(_4862_) );
AOI22X1 AOI22X1_282 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[346]), .C(w_mem_inst_w_mem_5__26_), .D(_4548__bF_buf5), .Y(_4863_) );
OAI21X1 OAI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_4862_), .B(_4547__bF_buf5), .C(_4863_), .Y(_3683__26_) );
AOI22X1 AOI22X1_283 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[347]), .C(w_mem_inst_w_mem_5__27_), .D(_4548__bF_buf4), .Y(_4864_) );
OAI21X1 OAI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_4406_), .B(_4547__bF_buf4), .C(_4864_), .Y(_3683__27_) );
INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__28_), .Y(_4865_) );
AOI22X1 AOI22X1_284 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[348]), .C(w_mem_inst_w_mem_5__28_), .D(_4548__bF_buf3), .Y(_4866_) );
OAI21X1 OAI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_4865_), .B(_4547__bF_buf3), .C(_4866_), .Y(_3683__28_) );
AOI22X1 AOI22X1_285 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[349]), .C(w_mem_inst_w_mem_5__29_), .D(_4548__bF_buf2), .Y(_4867_) );
OAI21X1 OAI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_4456_), .B(_4547__bF_buf2), .C(_4867_), .Y(_3683__29_) );
INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__30_), .Y(_4868_) );
AOI22X1 AOI22X1_286 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[350]), .C(w_mem_inst_w_mem_5__30_), .D(_4548__bF_buf1), .Y(_4869_) );
OAI21X1 OAI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_4868_), .B(_4547__bF_buf1), .C(_4869_), .Y(_3683__30_) );
AOI22X1 AOI22X1_287 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[351]), .C(w_mem_inst_w_mem_5__31_), .D(_4548__bF_buf0), .Y(_4870_) );
OAI21X1 OAI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_4509_), .B(_4547__bF_buf0), .C(_4870_), .Y(_3683__31_) );
INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__0_), .Y(_4871_) );
AOI22X1 AOI22X1_288 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[288]), .C(w_mem_inst_w_mem_6__0_), .D(_4548__bF_buf63), .Y(_4872_) );
OAI21X1 OAI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_4871_), .B(_4547__bF_buf63), .C(_4872_), .Y(_3684__0_) );
INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__1_), .Y(_4873_) );
AOI22X1 AOI22X1_289 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[289]), .C(w_mem_inst_w_mem_6__1_), .D(_4548__bF_buf62), .Y(_4874_) );
OAI21X1 OAI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_4873_), .B(_4547__bF_buf62), .C(_4874_), .Y(_3684__1_) );
INVX1 INVX1_264 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__2_), .Y(_4875_) );
AOI22X1 AOI22X1_290 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[290]), .C(w_mem_inst_w_mem_6__2_), .D(_4548__bF_buf61), .Y(_4876_) );
OAI21X1 OAI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_4875_), .B(_4547__bF_buf61), .C(_4876_), .Y(_3684__2_) );
INVX1 INVX1_265 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__3_), .Y(_4877_) );
AOI22X1 AOI22X1_291 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[291]), .C(w_mem_inst_w_mem_6__3_), .D(_4548__bF_buf60), .Y(_4878_) );
OAI21X1 OAI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_4877_), .B(_4547__bF_buf60), .C(_4878_), .Y(_3684__3_) );
AOI22X1 AOI22X1_292 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[292]), .C(w_mem_inst_w_mem_6__4_), .D(_4548__bF_buf59), .Y(_4879_) );
OAI21X1 OAI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3835_), .B(_4547__bF_buf59), .C(_4879_), .Y(_3684__4_) );
INVX1 INVX1_266 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__5_), .Y(_4880_) );
AOI22X1 AOI22X1_293 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[293]), .C(w_mem_inst_w_mem_6__5_), .D(_4548__bF_buf58), .Y(_4881_) );
OAI21X1 OAI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_4880_), .B(_4547__bF_buf58), .C(_4881_), .Y(_3684__5_) );
AOI22X1 AOI22X1_294 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[294]), .C(w_mem_inst_w_mem_6__6_), .D(_4548__bF_buf57), .Y(_4882_) );
OAI21X1 OAI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_3888_), .B(_4547__bF_buf57), .C(_4882_), .Y(_3684__6_) );
INVX1 INVX1_267 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__7_), .Y(_4883_) );
AOI22X1 AOI22X1_295 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[295]), .C(w_mem_inst_w_mem_6__7_), .D(_4548__bF_buf56), .Y(_4884_) );
OAI21X1 OAI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_4883_), .B(_4547__bF_buf56), .C(_4884_), .Y(_3684__7_) );
AOI22X1 AOI22X1_296 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[296]), .C(w_mem_inst_w_mem_6__8_), .D(_4548__bF_buf55), .Y(_4885_) );
OAI21X1 OAI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_3938_), .B(_4547__bF_buf55), .C(_4885_), .Y(_3684__8_) );
INVX1 INVX1_268 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__9_), .Y(_4886_) );
AOI22X1 AOI22X1_297 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[297]), .C(w_mem_inst_w_mem_6__9_), .D(_4548__bF_buf54), .Y(_4887_) );
OAI21X1 OAI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_4886_), .B(_4547__bF_buf54), .C(_4887_), .Y(_3684__9_) );
INVX1 INVX1_269 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__10_), .Y(_4888_) );
AOI22X1 AOI22X1_298 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[298]), .C(w_mem_inst_w_mem_6__10_), .D(_4548__bF_buf53), .Y(_4889_) );
OAI21X1 OAI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_4888_), .B(_4547__bF_buf53), .C(_4889_), .Y(_3684__10_) );
INVX1 INVX1_270 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__11_), .Y(_4890_) );
AOI22X1 AOI22X1_299 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[299]), .C(w_mem_inst_w_mem_6__11_), .D(_4548__bF_buf52), .Y(_4891_) );
OAI21X1 OAI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_4890_), .B(_4547__bF_buf52), .C(_4891_), .Y(_3684__11_) );
AOI22X1 AOI22X1_300 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[300]), .C(w_mem_inst_w_mem_6__12_), .D(_4548__bF_buf51), .Y(_4892_) );
OAI21X1 OAI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_4036_), .B(_4547__bF_buf51), .C(_4892_), .Y(_3684__12_) );
INVX1 INVX1_271 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__13_), .Y(_4893_) );
AOI22X1 AOI22X1_301 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[301]), .C(w_mem_inst_w_mem_6__13_), .D(_4548__bF_buf50), .Y(_4894_) );
OAI21X1 OAI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_4893_), .B(_4547__bF_buf50), .C(_4894_), .Y(_3684__13_) );
AOI22X1 AOI22X1_302 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[302]), .C(w_mem_inst_w_mem_6__14_), .D(_4548__bF_buf49), .Y(_4895_) );
OAI21X1 OAI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_4086_), .B(_4547__bF_buf49), .C(_4895_), .Y(_3684__14_) );
INVX1 INVX1_272 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__15_), .Y(_4896_) );
AOI22X1 AOI22X1_303 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[303]), .C(w_mem_inst_w_mem_6__15_), .D(_4548__bF_buf48), .Y(_4897_) );
OAI21X1 OAI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_4896_), .B(_4547__bF_buf48), .C(_4897_), .Y(_3684__15_) );
AOI22X1 AOI22X1_304 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[304]), .C(w_mem_inst_w_mem_6__16_), .D(_4548__bF_buf47), .Y(_4898_) );
OAI21X1 OAI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_4136_), .B(_4547__bF_buf47), .C(_4898_), .Y(_3684__16_) );
INVX1 INVX1_273 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__17_), .Y(_4899_) );
AOI22X1 AOI22X1_305 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[305]), .C(w_mem_inst_w_mem_6__17_), .D(_4548__bF_buf46), .Y(_4900_) );
OAI21X1 OAI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_4899_), .B(_4547__bF_buf46), .C(_4900_), .Y(_3684__17_) );
INVX1 INVX1_274 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__18_), .Y(_4901_) );
AOI22X1 AOI22X1_306 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[306]), .C(w_mem_inst_w_mem_6__18_), .D(_4548__bF_buf45), .Y(_4902_) );
OAI21X1 OAI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_4901_), .B(_4547__bF_buf45), .C(_4902_), .Y(_3684__18_) );
INVX1 INVX1_275 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__19_), .Y(_4903_) );
AOI22X1 AOI22X1_307 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[307]), .C(w_mem_inst_w_mem_6__19_), .D(_4548__bF_buf44), .Y(_4904_) );
OAI21X1 OAI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_4903_), .B(_4547__bF_buf44), .C(_4904_), .Y(_3684__19_) );
AOI22X1 AOI22X1_308 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[308]), .C(w_mem_inst_w_mem_6__20_), .D(_4548__bF_buf43), .Y(_4905_) );
OAI21X1 OAI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_4234_), .B(_4547__bF_buf43), .C(_4905_), .Y(_3684__20_) );
INVX1 INVX1_276 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__21_), .Y(_4906_) );
AOI22X1 AOI22X1_309 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[309]), .C(w_mem_inst_w_mem_6__21_), .D(_4548__bF_buf42), .Y(_4907_) );
OAI21X1 OAI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_4906_), .B(_4547__bF_buf42), .C(_4907_), .Y(_3684__21_) );
AOI22X1 AOI22X1_310 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[310]), .C(w_mem_inst_w_mem_6__22_), .D(_4548__bF_buf41), .Y(_4908_) );
OAI21X1 OAI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_4284_), .B(_4547__bF_buf41), .C(_4908_), .Y(_3684__22_) );
INVX1 INVX1_277 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__23_), .Y(_4909_) );
AOI22X1 AOI22X1_311 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[311]), .C(w_mem_inst_w_mem_6__23_), .D(_4548__bF_buf40), .Y(_4910_) );
OAI21X1 OAI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_4909_), .B(_4547__bF_buf40), .C(_4910_), .Y(_3684__23_) );
AOI22X1 AOI22X1_312 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[312]), .C(w_mem_inst_w_mem_6__24_), .D(_4548__bF_buf39), .Y(_4911_) );
OAI21X1 OAI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_4334_), .B(_4547__bF_buf39), .C(_4911_), .Y(_3684__24_) );
INVX1 INVX1_278 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__25_), .Y(_4912_) );
AOI22X1 AOI22X1_313 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[313]), .C(w_mem_inst_w_mem_6__25_), .D(_4548__bF_buf38), .Y(_4913_) );
OAI21X1 OAI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_4912_), .B(_4547__bF_buf38), .C(_4913_), .Y(_3684__25_) );
INVX1 INVX1_279 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__26_), .Y(_4914_) );
AOI22X1 AOI22X1_314 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[314]), .C(w_mem_inst_w_mem_6__26_), .D(_4548__bF_buf37), .Y(_4915_) );
OAI21X1 OAI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_4914_), .B(_4547__bF_buf37), .C(_4915_), .Y(_3684__26_) );
INVX1 INVX1_280 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__27_), .Y(_4916_) );
AOI22X1 AOI22X1_315 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[315]), .C(w_mem_inst_w_mem_6__27_), .D(_4548__bF_buf36), .Y(_4917_) );
OAI21X1 OAI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_4916_), .B(_4547__bF_buf36), .C(_4917_), .Y(_3684__27_) );
AOI22X1 AOI22X1_316 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[316]), .C(w_mem_inst_w_mem_6__28_), .D(_4548__bF_buf35), .Y(_4918_) );
OAI21X1 OAI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_4432_), .B(_4547__bF_buf35), .C(_4918_), .Y(_3684__28_) );
INVX1 INVX1_281 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__29_), .Y(_4919_) );
AOI22X1 AOI22X1_317 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[317]), .C(w_mem_inst_w_mem_6__29_), .D(_4548__bF_buf34), .Y(_4920_) );
OAI21X1 OAI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_4919_), .B(_4547__bF_buf34), .C(_4920_), .Y(_3684__29_) );
AOI22X1 AOI22X1_318 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[318]), .C(w_mem_inst_w_mem_6__30_), .D(_4548__bF_buf33), .Y(_4921_) );
OAI21X1 OAI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_4482_), .B(_4547__bF_buf33), .C(_4921_), .Y(_3684__30_) );
AOI22X1 AOI22X1_319 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[319]), .C(w_mem_inst_w_mem_6__31_), .D(_4548__bF_buf32), .Y(_4922_) );
OAI21X1 OAI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_4505_), .B(_4547__bF_buf32), .C(_4922_), .Y(_3684__31_) );
AOI22X1 AOI22X1_320 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[256]), .C(w_mem_inst_w_mem_7__0_), .D(_4548__bF_buf31), .Y(_4923_) );
OAI21X1 OAI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_3713_), .B(_4547__bF_buf31), .C(_4923_), .Y(_3685__0_) );
INVX1 INVX1_282 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__1_), .Y(_4924_) );
AOI22X1 AOI22X1_321 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[257]), .C(w_mem_inst_w_mem_7__1_), .D(_4548__bF_buf30), .Y(_4925_) );
OAI21X1 OAI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_4924_), .B(_4547__bF_buf30), .C(_4925_), .Y(_3685__1_) );
INVX1 INVX1_283 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__2_), .Y(_4926_) );
AOI22X1 AOI22X1_322 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[258]), .C(w_mem_inst_w_mem_7__2_), .D(_4548__bF_buf29), .Y(_4927_) );
OAI21X1 OAI21X1_285 ( .gnd(gnd), .vdd(vdd), .A(_4926_), .B(_4547__bF_buf29), .C(_4927_), .Y(_3685__2_) );
INVX1 INVX1_284 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__3_), .Y(_4928_) );
AOI22X1 AOI22X1_323 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[259]), .C(w_mem_inst_w_mem_7__3_), .D(_4548__bF_buf28), .Y(_4929_) );
OAI21X1 OAI21X1_286 ( .gnd(gnd), .vdd(vdd), .A(_4928_), .B(_4547__bF_buf28), .C(_4929_), .Y(_3685__3_) );
INVX1 INVX1_285 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__4_), .Y(_4930_) );
AOI22X1 AOI22X1_324 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[260]), .C(w_mem_inst_w_mem_7__4_), .D(_4548__bF_buf27), .Y(_4931_) );
OAI21X1 OAI21X1_287 ( .gnd(gnd), .vdd(vdd), .A(_4930_), .B(_4547__bF_buf27), .C(_4931_), .Y(_3685__4_) );
AOI22X1 AOI22X1_325 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[261]), .C(w_mem_inst_w_mem_7__5_), .D(_4548__bF_buf26), .Y(_4932_) );
OAI21X1 OAI21X1_288 ( .gnd(gnd), .vdd(vdd), .A(_3860_), .B(_4547__bF_buf26), .C(_4932_), .Y(_3685__5_) );
INVX1 INVX1_286 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__6_), .Y(_4933_) );
AOI22X1 AOI22X1_326 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[262]), .C(w_mem_inst_w_mem_7__6_), .D(_4548__bF_buf25), .Y(_4934_) );
OAI21X1 OAI21X1_289 ( .gnd(gnd), .vdd(vdd), .A(_4933_), .B(_4547__bF_buf25), .C(_4934_), .Y(_3685__6_) );
INVX1 INVX1_287 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__7_), .Y(_4935_) );
AOI22X1 AOI22X1_327 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[263]), .C(w_mem_inst_w_mem_7__7_), .D(_4548__bF_buf24), .Y(_4936_) );
OAI21X1 OAI21X1_290 ( .gnd(gnd), .vdd(vdd), .A(_4935_), .B(_4547__bF_buf24), .C(_4936_), .Y(_3685__7_) );
AOI22X1 AOI22X1_328 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[264]), .C(w_mem_inst_w_mem_7__8_), .D(_4548__bF_buf23), .Y(_4937_) );
OAI21X1 OAI21X1_291 ( .gnd(gnd), .vdd(vdd), .A(_3936_), .B(_4547__bF_buf23), .C(_4937_), .Y(_3685__8_) );
AOI22X1 AOI22X1_329 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[265]), .C(w_mem_inst_w_mem_7__9_), .D(_4548__bF_buf22), .Y(_4938_) );
OAI21X1 OAI21X1_292 ( .gnd(gnd), .vdd(vdd), .A(_3963_), .B(_4547__bF_buf22), .C(_4938_), .Y(_3685__9_) );
AOI22X1 AOI22X1_330 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[266]), .C(w_mem_inst_w_mem_7__10_), .D(_4548__bF_buf21), .Y(_4939_) );
OAI21X1 OAI21X1_293 ( .gnd(gnd), .vdd(vdd), .A(_3988_), .B(_4547__bF_buf21), .C(_4939_), .Y(_3685__10_) );
AOI22X1 AOI22X1_331 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[267]), .C(w_mem_inst_w_mem_7__11_), .D(_4548__bF_buf20), .Y(_4940_) );
OAI21X1 OAI21X1_294 ( .gnd(gnd), .vdd(vdd), .A(_4013_), .B(_4547__bF_buf20), .C(_4940_), .Y(_3685__11_) );
INVX1 INVX1_288 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__12_), .Y(_4941_) );
AOI22X1 AOI22X1_332 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[268]), .C(w_mem_inst_w_mem_7__12_), .D(_4548__bF_buf19), .Y(_4942_) );
OAI21X1 OAI21X1_295 ( .gnd(gnd), .vdd(vdd), .A(_4941_), .B(_4547__bF_buf19), .C(_4942_), .Y(_3685__12_) );
AOI22X1 AOI22X1_333 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[269]), .C(w_mem_inst_w_mem_7__13_), .D(_4548__bF_buf18), .Y(_4943_) );
OAI21X1 OAI21X1_296 ( .gnd(gnd), .vdd(vdd), .A(_4063_), .B(_4547__bF_buf18), .C(_4943_), .Y(_3685__13_) );
INVX1 INVX1_289 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__14_), .Y(_4944_) );
AOI22X1 AOI22X1_334 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[270]), .C(w_mem_inst_w_mem_7__14_), .D(_4548__bF_buf17), .Y(_4945_) );
OAI21X1 OAI21X1_297 ( .gnd(gnd), .vdd(vdd), .A(_4944_), .B(_4547__bF_buf17), .C(_4945_), .Y(_3685__14_) );
INVX1 INVX1_290 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__15_), .Y(_4946_) );
AOI22X1 AOI22X1_335 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[271]), .C(w_mem_inst_w_mem_7__15_), .D(_4548__bF_buf16), .Y(_4947_) );
OAI21X1 OAI21X1_298 ( .gnd(gnd), .vdd(vdd), .A(_4946_), .B(_4547__bF_buf16), .C(_4947_), .Y(_3685__15_) );
AOI22X1 AOI22X1_336 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[272]), .C(w_mem_inst_w_mem_7__16_), .D(_4548__bF_buf15), .Y(_4948_) );
OAI21X1 OAI21X1_299 ( .gnd(gnd), .vdd(vdd), .A(_4134_), .B(_4547__bF_buf15), .C(_4948_), .Y(_3685__16_) );
AOI22X1 AOI22X1_337 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[273]), .C(w_mem_inst_w_mem_7__17_), .D(_4548__bF_buf14), .Y(_4949_) );
OAI21X1 OAI21X1_300 ( .gnd(gnd), .vdd(vdd), .A(_4161_), .B(_4547__bF_buf14), .C(_4949_), .Y(_3685__17_) );
AOI22X1 AOI22X1_338 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[274]), .C(w_mem_inst_w_mem_7__18_), .D(_4548__bF_buf13), .Y(_4950_) );
OAI21X1 OAI21X1_301 ( .gnd(gnd), .vdd(vdd), .A(_4186_), .B(_4547__bF_buf13), .C(_4950_), .Y(_3685__18_) );
AOI22X1 AOI22X1_339 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[275]), .C(w_mem_inst_w_mem_7__19_), .D(_4548__bF_buf12), .Y(_4951_) );
OAI21X1 OAI21X1_302 ( .gnd(gnd), .vdd(vdd), .A(_4211_), .B(_4547__bF_buf12), .C(_4951_), .Y(_3685__19_) );
INVX1 INVX1_291 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__20_), .Y(_4952_) );
AOI22X1 AOI22X1_340 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[276]), .C(w_mem_inst_w_mem_7__20_), .D(_4548__bF_buf11), .Y(_4953_) );
OAI21X1 OAI21X1_303 ( .gnd(gnd), .vdd(vdd), .A(_4952_), .B(_4547__bF_buf11), .C(_4953_), .Y(_3685__20_) );
AOI22X1 AOI22X1_341 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[277]), .C(w_mem_inst_w_mem_7__21_), .D(_4548__bF_buf10), .Y(_4954_) );
OAI21X1 OAI21X1_304 ( .gnd(gnd), .vdd(vdd), .A(_4261_), .B(_4547__bF_buf10), .C(_4954_), .Y(_3685__21_) );
INVX1 INVX1_292 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__22_), .Y(_4955_) );
AOI22X1 AOI22X1_342 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[278]), .C(w_mem_inst_w_mem_7__22_), .D(_4548__bF_buf9), .Y(_4956_) );
OAI21X1 OAI21X1_305 ( .gnd(gnd), .vdd(vdd), .A(_4955_), .B(_4547__bF_buf9), .C(_4956_), .Y(_3685__22_) );
INVX1 INVX1_293 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__23_), .Y(_4957_) );
AOI22X1 AOI22X1_343 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[279]), .C(w_mem_inst_w_mem_7__23_), .D(_4548__bF_buf8), .Y(_4958_) );
OAI21X1 OAI21X1_306 ( .gnd(gnd), .vdd(vdd), .A(_4957_), .B(_4547__bF_buf8), .C(_4958_), .Y(_3685__23_) );
AOI22X1 AOI22X1_344 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[280]), .C(w_mem_inst_w_mem_7__24_), .D(_4548__bF_buf7), .Y(_4959_) );
OAI21X1 OAI21X1_307 ( .gnd(gnd), .vdd(vdd), .A(_4332_), .B(_4547__bF_buf7), .C(_4959_), .Y(_3685__24_) );
AOI22X1 AOI22X1_345 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[281]), .C(w_mem_inst_w_mem_7__25_), .D(_4548__bF_buf6), .Y(_4960_) );
OAI21X1 OAI21X1_308 ( .gnd(gnd), .vdd(vdd), .A(_4359_), .B(_4547__bF_buf6), .C(_4960_), .Y(_3685__25_) );
AOI22X1 AOI22X1_346 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[282]), .C(w_mem_inst_w_mem_7__26_), .D(_4548__bF_buf5), .Y(_4961_) );
OAI21X1 OAI21X1_309 ( .gnd(gnd), .vdd(vdd), .A(_4384_), .B(_4547__bF_buf5), .C(_4961_), .Y(_3685__26_) );
AOI22X1 AOI22X1_347 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[283]), .C(w_mem_inst_w_mem_7__27_), .D(_4548__bF_buf4), .Y(_4962_) );
OAI21X1 OAI21X1_310 ( .gnd(gnd), .vdd(vdd), .A(_4409_), .B(_4547__bF_buf4), .C(_4962_), .Y(_3685__27_) );
INVX1 INVX1_294 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__28_), .Y(_4963_) );
AOI22X1 AOI22X1_348 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[284]), .C(w_mem_inst_w_mem_7__28_), .D(_4548__bF_buf3), .Y(_4964_) );
OAI21X1 OAI21X1_311 ( .gnd(gnd), .vdd(vdd), .A(_4963_), .B(_4547__bF_buf3), .C(_4964_), .Y(_3685__28_) );
AOI22X1 AOI22X1_349 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[285]), .C(w_mem_inst_w_mem_7__29_), .D(_4548__bF_buf2), .Y(_4965_) );
OAI21X1 OAI21X1_312 ( .gnd(gnd), .vdd(vdd), .A(_4459_), .B(_4547__bF_buf2), .C(_4965_), .Y(_3685__29_) );
INVX1 INVX1_295 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__30_), .Y(_4966_) );
AOI22X1 AOI22X1_350 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[286]), .C(w_mem_inst_w_mem_7__30_), .D(_4548__bF_buf1), .Y(_4967_) );
OAI21X1 OAI21X1_313 ( .gnd(gnd), .vdd(vdd), .A(_4966_), .B(_4547__bF_buf1), .C(_4967_), .Y(_3685__30_) );
INVX1 INVX1_296 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__31_), .Y(_4968_) );
AOI22X1 AOI22X1_351 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[287]), .C(w_mem_inst_w_mem_7__31_), .D(_4548__bF_buf0), .Y(_4969_) );
OAI21X1 OAI21X1_314 ( .gnd(gnd), .vdd(vdd), .A(_4968_), .B(_4547__bF_buf0), .C(_4969_), .Y(_3685__31_) );
INVX1 INVX1_297 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__0_), .Y(_4970_) );
AOI22X1 AOI22X1_352 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[224]), .C(w_mem_inst_w_mem_8__0_), .D(_4548__bF_buf63), .Y(_4971_) );
OAI21X1 OAI21X1_315 ( .gnd(gnd), .vdd(vdd), .A(_4970_), .B(_4547__bF_buf63), .C(_4971_), .Y(_3686__0_) );
AOI22X1 AOI22X1_353 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[225]), .C(w_mem_inst_w_mem_8__1_), .D(_4548__bF_buf62), .Y(_4972_) );
OAI21X1 OAI21X1_316 ( .gnd(gnd), .vdd(vdd), .A(_3761_), .B(_4547__bF_buf62), .C(_4972_), .Y(_3686__1_) );
AOI22X1 AOI22X1_354 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[226]), .C(w_mem_inst_w_mem_8__2_), .D(_4548__bF_buf61), .Y(_4973_) );
OAI21X1 OAI21X1_317 ( .gnd(gnd), .vdd(vdd), .A(_3785_), .B(_4547__bF_buf61), .C(_4973_), .Y(_3686__2_) );
AOI22X1 AOI22X1_355 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[227]), .C(w_mem_inst_w_mem_8__3_), .D(_4548__bF_buf60), .Y(_4974_) );
OAI21X1 OAI21X1_318 ( .gnd(gnd), .vdd(vdd), .A(_3813_), .B(_4547__bF_buf60), .C(_4974_), .Y(_3686__3_) );
AOI22X1 AOI22X1_356 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[228]), .C(w_mem_inst_w_mem_8__4_), .D(_4548__bF_buf59), .Y(_4975_) );
OAI21X1 OAI21X1_319 ( .gnd(gnd), .vdd(vdd), .A(_3840_), .B(_4547__bF_buf59), .C(_4975_), .Y(_3686__4_) );
AOI22X1 AOI22X1_357 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[229]), .C(w_mem_inst_w_mem_8__5_), .D(_4548__bF_buf58), .Y(_4976_) );
OAI21X1 OAI21X1_320 ( .gnd(gnd), .vdd(vdd), .A(_3862_), .B(_4547__bF_buf58), .C(_4976_), .Y(_3686__5_) );
AOI22X1 AOI22X1_358 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[230]), .C(w_mem_inst_w_mem_8__6_), .D(_4548__bF_buf57), .Y(_4977_) );
OAI21X1 OAI21X1_321 ( .gnd(gnd), .vdd(vdd), .A(_3887_), .B(_4547__bF_buf57), .C(_4977_), .Y(_3686__6_) );
INVX1 INVX1_298 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__7_), .Y(_4978_) );
AOI22X1 AOI22X1_359 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[231]), .C(w_mem_inst_w_mem_8__7_), .D(_4548__bF_buf56), .Y(_4979_) );
OAI21X1 OAI21X1_322 ( .gnd(gnd), .vdd(vdd), .A(_4978_), .B(_4547__bF_buf56), .C(_4979_), .Y(_3686__7_) );
INVX1 INVX1_299 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__8_), .Y(_4980_) );
AOI22X1 AOI22X1_360 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[232]), .C(w_mem_inst_w_mem_8__8_), .D(_4548__bF_buf55), .Y(_4981_) );
OAI21X1 OAI21X1_323 ( .gnd(gnd), .vdd(vdd), .A(_4980_), .B(_4547__bF_buf55), .C(_4981_), .Y(_3686__8_) );
INVX1 INVX1_300 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__9_), .Y(_4982_) );
AOI22X1 AOI22X1_361 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[233]), .C(w_mem_inst_w_mem_8__9_), .D(_4548__bF_buf54), .Y(_4983_) );
OAI21X1 OAI21X1_324 ( .gnd(gnd), .vdd(vdd), .A(_4982_), .B(_4547__bF_buf54), .C(_4983_), .Y(_3686__9_) );
INVX1 INVX1_301 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__10_), .Y(_4984_) );
AOI22X1 AOI22X1_362 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[234]), .C(w_mem_inst_w_mem_8__10_), .D(_4548__bF_buf53), .Y(_4985_) );
OAI21X1 OAI21X1_325 ( .gnd(gnd), .vdd(vdd), .A(_4984_), .B(_4547__bF_buf53), .C(_4985_), .Y(_3686__10_) );
INVX1 INVX1_302 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__11_), .Y(_4986_) );
AOI22X1 AOI22X1_363 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[235]), .C(w_mem_inst_w_mem_8__11_), .D(_4548__bF_buf52), .Y(_4987_) );
OAI21X1 OAI21X1_326 ( .gnd(gnd), .vdd(vdd), .A(_4986_), .B(_4547__bF_buf52), .C(_4987_), .Y(_3686__11_) );
AOI22X1 AOI22X1_364 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[236]), .C(w_mem_inst_w_mem_8__12_), .D(_4548__bF_buf51), .Y(_4988_) );
OAI21X1 OAI21X1_327 ( .gnd(gnd), .vdd(vdd), .A(_4035_), .B(_4547__bF_buf51), .C(_4988_), .Y(_3686__12_) );
INVX1 INVX1_303 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__13_), .Y(_4989_) );
AOI22X1 AOI22X1_365 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[237]), .C(w_mem_inst_w_mem_8__13_), .D(_4548__bF_buf50), .Y(_4990_) );
OAI21X1 OAI21X1_328 ( .gnd(gnd), .vdd(vdd), .A(_4989_), .B(_4547__bF_buf50), .C(_4990_), .Y(_3686__13_) );
AOI22X1 AOI22X1_366 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[238]), .C(w_mem_inst_w_mem_8__14_), .D(_4548__bF_buf49), .Y(_4991_) );
OAI21X1 OAI21X1_329 ( .gnd(gnd), .vdd(vdd), .A(_4085_), .B(_4547__bF_buf49), .C(_4991_), .Y(_3686__14_) );
INVX1 INVX1_304 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__15_), .Y(_4992_) );
AOI22X1 AOI22X1_367 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[239]), .C(w_mem_inst_w_mem_8__15_), .D(_4548__bF_buf48), .Y(_4993_) );
OAI21X1 OAI21X1_330 ( .gnd(gnd), .vdd(vdd), .A(_4992_), .B(_4547__bF_buf48), .C(_4993_), .Y(_3686__15_) );
INVX1 INVX1_305 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__16_), .Y(_4994_) );
AOI22X1 AOI22X1_368 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[240]), .C(w_mem_inst_w_mem_8__16_), .D(_4548__bF_buf47), .Y(_4995_) );
OAI21X1 OAI21X1_331 ( .gnd(gnd), .vdd(vdd), .A(_4994_), .B(_4547__bF_buf47), .C(_4995_), .Y(_3686__16_) );
INVX1 INVX1_306 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__17_), .Y(_4996_) );
AOI22X1 AOI22X1_369 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[241]), .C(w_mem_inst_w_mem_8__17_), .D(_4548__bF_buf46), .Y(_4997_) );
OAI21X1 OAI21X1_332 ( .gnd(gnd), .vdd(vdd), .A(_4996_), .B(_4547__bF_buf46), .C(_4997_), .Y(_3686__17_) );
INVX1 INVX1_307 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__18_), .Y(_4998_) );
AOI22X1 AOI22X1_370 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[242]), .C(w_mem_inst_w_mem_8__18_), .D(_4548__bF_buf45), .Y(_4999_) );
OAI21X1 OAI21X1_333 ( .gnd(gnd), .vdd(vdd), .A(_4998_), .B(_4547__bF_buf45), .C(_4999_), .Y(_3686__18_) );
INVX1 INVX1_308 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__19_), .Y(_5000_) );
AOI22X1 AOI22X1_371 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[243]), .C(w_mem_inst_w_mem_8__19_), .D(_4548__bF_buf44), .Y(_5001_) );
OAI21X1 OAI21X1_334 ( .gnd(gnd), .vdd(vdd), .A(_5000_), .B(_4547__bF_buf44), .C(_5001_), .Y(_3686__19_) );
AOI22X1 AOI22X1_372 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[244]), .C(w_mem_inst_w_mem_8__20_), .D(_4548__bF_buf43), .Y(_5002_) );
OAI21X1 OAI21X1_335 ( .gnd(gnd), .vdd(vdd), .A(_4233_), .B(_4547__bF_buf43), .C(_5002_), .Y(_3686__20_) );
INVX1 INVX1_309 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__21_), .Y(_5003_) );
AOI22X1 AOI22X1_373 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[245]), .C(w_mem_inst_w_mem_8__21_), .D(_4548__bF_buf42), .Y(_5004_) );
OAI21X1 OAI21X1_336 ( .gnd(gnd), .vdd(vdd), .A(_5003_), .B(_4547__bF_buf42), .C(_5004_), .Y(_3686__21_) );
AOI22X1 AOI22X1_374 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[246]), .C(w_mem_inst_w_mem_8__22_), .D(_4548__bF_buf41), .Y(_5005_) );
OAI21X1 OAI21X1_337 ( .gnd(gnd), .vdd(vdd), .A(_4283_), .B(_4547__bF_buf41), .C(_5005_), .Y(_3686__22_) );
INVX1 INVX1_310 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__23_), .Y(_5006_) );
AOI22X1 AOI22X1_375 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[247]), .C(w_mem_inst_w_mem_8__23_), .D(_4548__bF_buf40), .Y(_5007_) );
OAI21X1 OAI21X1_338 ( .gnd(gnd), .vdd(vdd), .A(_5006_), .B(_4547__bF_buf40), .C(_5007_), .Y(_3686__23_) );
INVX1 INVX1_311 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__24_), .Y(_5008_) );
AOI22X1 AOI22X1_376 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[248]), .C(w_mem_inst_w_mem_8__24_), .D(_4548__bF_buf39), .Y(_5009_) );
OAI21X1 OAI21X1_339 ( .gnd(gnd), .vdd(vdd), .A(_5008_), .B(_4547__bF_buf39), .C(_5009_), .Y(_3686__24_) );
INVX1 INVX1_312 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__25_), .Y(_5010_) );
AOI22X1 AOI22X1_377 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[249]), .C(w_mem_inst_w_mem_8__25_), .D(_4548__bF_buf38), .Y(_5011_) );
OAI21X1 OAI21X1_340 ( .gnd(gnd), .vdd(vdd), .A(_5010_), .B(_4547__bF_buf38), .C(_5011_), .Y(_3686__25_) );
INVX1 INVX1_313 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__26_), .Y(_5012_) );
AOI22X1 AOI22X1_378 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[250]), .C(w_mem_inst_w_mem_8__26_), .D(_4548__bF_buf37), .Y(_5013_) );
OAI21X1 OAI21X1_341 ( .gnd(gnd), .vdd(vdd), .A(_5012_), .B(_4547__bF_buf37), .C(_5013_), .Y(_3686__26_) );
INVX1 INVX1_314 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__27_), .Y(_5014_) );
AOI22X1 AOI22X1_379 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[251]), .C(w_mem_inst_w_mem_8__27_), .D(_4548__bF_buf36), .Y(_5015_) );
OAI21X1 OAI21X1_342 ( .gnd(gnd), .vdd(vdd), .A(_5014_), .B(_4547__bF_buf36), .C(_5015_), .Y(_3686__27_) );
AOI22X1 AOI22X1_380 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[252]), .C(w_mem_inst_w_mem_8__28_), .D(_4548__bF_buf35), .Y(_5016_) );
OAI21X1 OAI21X1_343 ( .gnd(gnd), .vdd(vdd), .A(_4431_), .B(_4547__bF_buf35), .C(_5016_), .Y(_3686__28_) );
INVX1 INVX1_315 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__29_), .Y(_5017_) );
AOI22X1 AOI22X1_381 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[253]), .C(w_mem_inst_w_mem_8__29_), .D(_4548__bF_buf34), .Y(_5018_) );
OAI21X1 OAI21X1_344 ( .gnd(gnd), .vdd(vdd), .A(_5017_), .B(_4547__bF_buf34), .C(_5018_), .Y(_3686__29_) );
AOI22X1 AOI22X1_382 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[254]), .C(w_mem_inst_w_mem_8__30_), .D(_4548__bF_buf33), .Y(_5019_) );
OAI21X1 OAI21X1_345 ( .gnd(gnd), .vdd(vdd), .A(_4481_), .B(_4547__bF_buf33), .C(_5019_), .Y(_3686__30_) );
AOI22X1 AOI22X1_383 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[255]), .C(w_mem_inst_w_mem_8__31_), .D(_4548__bF_buf32), .Y(_5020_) );
OAI21X1 OAI21X1_346 ( .gnd(gnd), .vdd(vdd), .A(_4508_), .B(_4547__bF_buf32), .C(_5020_), .Y(_3686__31_) );
INVX1 INVX1_316 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__0_), .Y(_5021_) );
AOI22X1 AOI22X1_384 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[192]), .C(w_mem_inst_w_mem_9__0_), .D(_4548__bF_buf31), .Y(_5022_) );
OAI21X1 OAI21X1_347 ( .gnd(gnd), .vdd(vdd), .A(_5021_), .B(_4547__bF_buf31), .C(_5022_), .Y(_3687__0_) );
INVX1 INVX1_317 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__1_), .Y(_5023_) );
AOI22X1 AOI22X1_385 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[193]), .C(w_mem_inst_w_mem_9__1_), .D(_4548__bF_buf30), .Y(_5024_) );
OAI21X1 OAI21X1_348 ( .gnd(gnd), .vdd(vdd), .A(_5023_), .B(_4547__bF_buf30), .C(_5024_), .Y(_3687__1_) );
AOI22X1 AOI22X1_386 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[194]), .C(w_mem_inst_w_mem_9__2_), .D(_4548__bF_buf29), .Y(_5025_) );
OAI21X1 OAI21X1_349 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(_4547__bF_buf29), .C(_5025_), .Y(_3687__2_) );
AOI22X1 AOI22X1_387 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[195]), .C(w_mem_inst_w_mem_9__3_), .D(_4548__bF_buf28), .Y(_5026_) );
OAI21X1 OAI21X1_350 ( .gnd(gnd), .vdd(vdd), .A(_3808_), .B(_4547__bF_buf28), .C(_5026_), .Y(_3687__3_) );
INVX1 INVX1_318 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__4_), .Y(_5027_) );
AOI22X1 AOI22X1_388 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[196]), .C(w_mem_inst_w_mem_9__4_), .D(_4548__bF_buf27), .Y(_5028_) );
OAI21X1 OAI21X1_351 ( .gnd(gnd), .vdd(vdd), .A(_5027_), .B(_4547__bF_buf27), .C(_5028_), .Y(_3687__4_) );
INVX1 INVX1_319 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__5_), .Y(_5029_) );
AOI22X1 AOI22X1_389 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[197]), .C(w_mem_inst_w_mem_9__5_), .D(_4548__bF_buf26), .Y(_5030_) );
OAI21X1 OAI21X1_352 ( .gnd(gnd), .vdd(vdd), .A(_5029_), .B(_4547__bF_buf26), .C(_5030_), .Y(_3687__5_) );
INVX1 INVX1_320 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__6_), .Y(_5031_) );
AOI22X1 AOI22X1_390 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[198]), .C(w_mem_inst_w_mem_9__6_), .D(_4548__bF_buf25), .Y(_5032_) );
OAI21X1 OAI21X1_353 ( .gnd(gnd), .vdd(vdd), .A(_5031_), .B(_4547__bF_buf25), .C(_5032_), .Y(_3687__6_) );
INVX1 INVX1_321 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__7_), .Y(_5033_) );
AOI22X1 AOI22X1_391 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[199]), .C(w_mem_inst_w_mem_9__7_), .D(_4548__bF_buf24), .Y(_5034_) );
OAI21X1 OAI21X1_354 ( .gnd(gnd), .vdd(vdd), .A(_5033_), .B(_4547__bF_buf24), .C(_5034_), .Y(_3687__7_) );
AOI22X1 AOI22X1_392 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[200]), .C(w_mem_inst_w_mem_9__8_), .D(_4548__bF_buf23), .Y(_5035_) );
OAI21X1 OAI21X1_355 ( .gnd(gnd), .vdd(vdd), .A(_3935_), .B(_4547__bF_buf23), .C(_5035_), .Y(_3687__8_) );
INVX1 INVX1_322 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__9_), .Y(_5036_) );
AOI22X1 AOI22X1_393 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[201]), .C(w_mem_inst_w_mem_9__9_), .D(_4548__bF_buf22), .Y(_5037_) );
OAI21X1 OAI21X1_356 ( .gnd(gnd), .vdd(vdd), .A(_5036_), .B(_4547__bF_buf22), .C(_5037_), .Y(_3687__9_) );
INVX1 INVX1_323 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__10_), .Y(_5038_) );
AOI22X1 AOI22X1_394 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[202]), .C(w_mem_inst_w_mem_9__10_), .D(_4548__bF_buf21), .Y(_5039_) );
OAI21X1 OAI21X1_357 ( .gnd(gnd), .vdd(vdd), .A(_5038_), .B(_4547__bF_buf21), .C(_5039_), .Y(_3687__10_) );
INVX1 INVX1_324 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__11_), .Y(_5040_) );
AOI22X1 AOI22X1_395 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[203]), .C(w_mem_inst_w_mem_9__11_), .D(_4548__bF_buf20), .Y(_5041_) );
OAI21X1 OAI21X1_358 ( .gnd(gnd), .vdd(vdd), .A(_5040_), .B(_4547__bF_buf20), .C(_5041_), .Y(_3687__11_) );
INVX1 INVX1_325 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__12_), .Y(_5042_) );
AOI22X1 AOI22X1_396 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[204]), .C(w_mem_inst_w_mem_9__12_), .D(_4548__bF_buf19), .Y(_5043_) );
OAI21X1 OAI21X1_359 ( .gnd(gnd), .vdd(vdd), .A(_5042_), .B(_4547__bF_buf19), .C(_5043_), .Y(_3687__12_) );
INVX1 INVX1_326 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__13_), .Y(_5044_) );
AOI22X1 AOI22X1_397 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[205]), .C(w_mem_inst_w_mem_9__13_), .D(_4548__bF_buf18), .Y(_5045_) );
OAI21X1 OAI21X1_360 ( .gnd(gnd), .vdd(vdd), .A(_5044_), .B(_4547__bF_buf18), .C(_5045_), .Y(_3687__13_) );
INVX1 INVX1_327 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__14_), .Y(_5046_) );
AOI22X1 AOI22X1_398 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[206]), .C(w_mem_inst_w_mem_9__14_), .D(_4548__bF_buf17), .Y(_5047_) );
OAI21X1 OAI21X1_361 ( .gnd(gnd), .vdd(vdd), .A(_5046_), .B(_4547__bF_buf17), .C(_5047_), .Y(_3687__14_) );
INVX1 INVX1_328 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__15_), .Y(_5048_) );
AOI22X1 AOI22X1_399 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[207]), .C(w_mem_inst_w_mem_9__15_), .D(_4548__bF_buf16), .Y(_5049_) );
OAI21X1 OAI21X1_362 ( .gnd(gnd), .vdd(vdd), .A(_5048_), .B(_4547__bF_buf16), .C(_5049_), .Y(_3687__15_) );
AOI22X1 AOI22X1_400 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[208]), .C(w_mem_inst_w_mem_9__16_), .D(_4548__bF_buf15), .Y(_5050_) );
OAI21X1 OAI21X1_363 ( .gnd(gnd), .vdd(vdd), .A(_4133_), .B(_4547__bF_buf15), .C(_5050_), .Y(_3687__16_) );
INVX1 INVX1_329 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__17_), .Y(_5051_) );
AOI22X1 AOI22X1_401 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[209]), .C(w_mem_inst_w_mem_9__17_), .D(_4548__bF_buf14), .Y(_5052_) );
OAI21X1 OAI21X1_364 ( .gnd(gnd), .vdd(vdd), .A(_5051_), .B(_4547__bF_buf14), .C(_5052_), .Y(_3687__17_) );
INVX1 INVX1_330 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__18_), .Y(_5053_) );
AOI22X1 AOI22X1_402 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[210]), .C(w_mem_inst_w_mem_9__18_), .D(_4548__bF_buf13), .Y(_5054_) );
OAI21X1 OAI21X1_365 ( .gnd(gnd), .vdd(vdd), .A(_5053_), .B(_4547__bF_buf13), .C(_5054_), .Y(_3687__18_) );
INVX1 INVX1_331 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__19_), .Y(_5055_) );
AOI22X1 AOI22X1_403 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[211]), .C(w_mem_inst_w_mem_9__19_), .D(_4548__bF_buf12), .Y(_5056_) );
OAI21X1 OAI21X1_366 ( .gnd(gnd), .vdd(vdd), .A(_5055_), .B(_4547__bF_buf12), .C(_5056_), .Y(_3687__19_) );
INVX1 INVX1_332 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__20_), .Y(_5057_) );
AOI22X1 AOI22X1_404 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[212]), .C(w_mem_inst_w_mem_9__20_), .D(_4548__bF_buf11), .Y(_5058_) );
OAI21X1 OAI21X1_367 ( .gnd(gnd), .vdd(vdd), .A(_5057_), .B(_4547__bF_buf11), .C(_5058_), .Y(_3687__20_) );
INVX1 INVX1_333 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__21_), .Y(_5059_) );
AOI22X1 AOI22X1_405 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[213]), .C(w_mem_inst_w_mem_9__21_), .D(_4548__bF_buf10), .Y(_5060_) );
OAI21X1 OAI21X1_368 ( .gnd(gnd), .vdd(vdd), .A(_5059_), .B(_4547__bF_buf10), .C(_5060_), .Y(_3687__21_) );
INVX1 INVX1_334 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__22_), .Y(_5061_) );
AOI22X1 AOI22X1_406 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[214]), .C(w_mem_inst_w_mem_9__22_), .D(_4548__bF_buf9), .Y(_5062_) );
OAI21X1 OAI21X1_369 ( .gnd(gnd), .vdd(vdd), .A(_5061_), .B(_4547__bF_buf9), .C(_5062_), .Y(_3687__22_) );
INVX1 INVX1_335 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__23_), .Y(_5063_) );
AOI22X1 AOI22X1_407 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[215]), .C(w_mem_inst_w_mem_9__23_), .D(_4548__bF_buf8), .Y(_5064_) );
OAI21X1 OAI21X1_370 ( .gnd(gnd), .vdd(vdd), .A(_5063_), .B(_4547__bF_buf8), .C(_5064_), .Y(_3687__23_) );
AOI22X1 AOI22X1_408 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[216]), .C(w_mem_inst_w_mem_9__24_), .D(_4548__bF_buf7), .Y(_5065_) );
OAI21X1 OAI21X1_371 ( .gnd(gnd), .vdd(vdd), .A(_4331_), .B(_4547__bF_buf7), .C(_5065_), .Y(_3687__24_) );
INVX1 INVX1_336 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__25_), .Y(_5066_) );
AOI22X1 AOI22X1_409 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[217]), .C(w_mem_inst_w_mem_9__25_), .D(_4548__bF_buf6), .Y(_5067_) );
OAI21X1 OAI21X1_372 ( .gnd(gnd), .vdd(vdd), .A(_5066_), .B(_4547__bF_buf6), .C(_5067_), .Y(_3687__25_) );
INVX1 INVX1_337 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__26_), .Y(_5068_) );
AOI22X1 AOI22X1_410 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[218]), .C(w_mem_inst_w_mem_9__26_), .D(_4548__bF_buf5), .Y(_5069_) );
OAI21X1 OAI21X1_373 ( .gnd(gnd), .vdd(vdd), .A(_5068_), .B(_4547__bF_buf5), .C(_5069_), .Y(_3687__26_) );
INVX1 INVX1_338 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__27_), .Y(_5070_) );
AOI22X1 AOI22X1_411 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[219]), .C(w_mem_inst_w_mem_9__27_), .D(_4548__bF_buf4), .Y(_5071_) );
OAI21X1 OAI21X1_374 ( .gnd(gnd), .vdd(vdd), .A(_5070_), .B(_4547__bF_buf4), .C(_5071_), .Y(_3687__27_) );
INVX1 INVX1_339 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__28_), .Y(_5072_) );
AOI22X1 AOI22X1_412 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[220]), .C(w_mem_inst_w_mem_9__28_), .D(_4548__bF_buf3), .Y(_5073_) );
OAI21X1 OAI21X1_375 ( .gnd(gnd), .vdd(vdd), .A(_5072_), .B(_4547__bF_buf3), .C(_5073_), .Y(_3687__28_) );
INVX1 INVX1_340 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__29_), .Y(_5074_) );
AOI22X1 AOI22X1_413 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[221]), .C(w_mem_inst_w_mem_9__29_), .D(_4548__bF_buf2), .Y(_5075_) );
OAI21X1 OAI21X1_376 ( .gnd(gnd), .vdd(vdd), .A(_5074_), .B(_4547__bF_buf2), .C(_5075_), .Y(_3687__29_) );
INVX1 INVX1_341 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__30_), .Y(_5076_) );
AOI22X1 AOI22X1_414 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[222]), .C(w_mem_inst_w_mem_9__30_), .D(_4548__bF_buf1), .Y(_5077_) );
OAI21X1 OAI21X1_377 ( .gnd(gnd), .vdd(vdd), .A(_5076_), .B(_4547__bF_buf1), .C(_5077_), .Y(_3687__30_) );
INVX1 INVX1_342 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__31_), .Y(_5078_) );
AOI22X1 AOI22X1_415 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[223]), .C(w_mem_inst_w_mem_9__31_), .D(_4548__bF_buf0), .Y(_5079_) );
OAI21X1 OAI21X1_378 ( .gnd(gnd), .vdd(vdd), .A(_5078_), .B(_4547__bF_buf0), .C(_5079_), .Y(_3687__31_) );
INVX1 INVX1_343 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__0_), .Y(_5080_) );
AOI22X1 AOI22X1_416 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[160]), .C(w_mem_inst_w_mem_10__0_), .D(_4548__bF_buf63), .Y(_5081_) );
OAI21X1 OAI21X1_379 ( .gnd(gnd), .vdd(vdd), .A(_5080_), .B(_4547__bF_buf63), .C(_5081_), .Y(_3673__0_) );
INVX1 INVX1_344 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__1_), .Y(_5082_) );
AOI22X1 AOI22X1_417 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[161]), .C(w_mem_inst_w_mem_10__1_), .D(_4548__bF_buf62), .Y(_5083_) );
OAI21X1 OAI21X1_380 ( .gnd(gnd), .vdd(vdd), .A(_5082_), .B(_4547__bF_buf62), .C(_5083_), .Y(_3673__1_) );
INVX1 INVX1_345 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__2_), .Y(_5084_) );
AOI22X1 AOI22X1_418 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[162]), .C(w_mem_inst_w_mem_10__2_), .D(_4548__bF_buf61), .Y(_5085_) );
OAI21X1 OAI21X1_381 ( .gnd(gnd), .vdd(vdd), .A(_5084_), .B(_4547__bF_buf61), .C(_5085_), .Y(_3673__2_) );
INVX1 INVX1_346 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__3_), .Y(_5086_) );
AOI22X1 AOI22X1_419 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[163]), .C(w_mem_inst_w_mem_10__3_), .D(_4548__bF_buf60), .Y(_5087_) );
OAI21X1 OAI21X1_382 ( .gnd(gnd), .vdd(vdd), .A(_5086_), .B(_4547__bF_buf60), .C(_5087_), .Y(_3673__3_) );
INVX1 INVX1_347 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__4_), .Y(_5088_) );
AOI22X1 AOI22X1_420 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[164]), .C(w_mem_inst_w_mem_10__4_), .D(_4548__bF_buf59), .Y(_5089_) );
OAI21X1 OAI21X1_383 ( .gnd(gnd), .vdd(vdd), .A(_5088_), .B(_4547__bF_buf59), .C(_5089_), .Y(_3673__4_) );
INVX1 INVX1_348 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__5_), .Y(_5090_) );
AOI22X1 AOI22X1_421 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[165]), .C(w_mem_inst_w_mem_10__5_), .D(_4548__bF_buf58), .Y(_5091_) );
OAI21X1 OAI21X1_384 ( .gnd(gnd), .vdd(vdd), .A(_5090_), .B(_4547__bF_buf58), .C(_5091_), .Y(_3673__5_) );
INVX1 INVX1_349 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__6_), .Y(_5092_) );
AOI22X1 AOI22X1_422 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[166]), .C(w_mem_inst_w_mem_10__6_), .D(_4548__bF_buf57), .Y(_5093_) );
OAI21X1 OAI21X1_385 ( .gnd(gnd), .vdd(vdd), .A(_5092_), .B(_4547__bF_buf57), .C(_5093_), .Y(_3673__6_) );
INVX1 INVX1_350 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__7_), .Y(_5094_) );
AOI22X1 AOI22X1_423 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[167]), .C(w_mem_inst_w_mem_10__7_), .D(_4548__bF_buf56), .Y(_5095_) );
OAI21X1 OAI21X1_386 ( .gnd(gnd), .vdd(vdd), .A(_5094_), .B(_4547__bF_buf56), .C(_5095_), .Y(_3673__7_) );
INVX1 INVX1_351 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__8_), .Y(_5096_) );
AOI22X1 AOI22X1_424 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[168]), .C(w_mem_inst_w_mem_10__8_), .D(_4548__bF_buf55), .Y(_5097_) );
OAI21X1 OAI21X1_387 ( .gnd(gnd), .vdd(vdd), .A(_5096_), .B(_4547__bF_buf55), .C(_5097_), .Y(_3673__8_) );
INVX1 INVX1_352 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__9_), .Y(_5098_) );
AOI22X1 AOI22X1_425 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[169]), .C(w_mem_inst_w_mem_10__9_), .D(_4548__bF_buf54), .Y(_5099_) );
OAI21X1 OAI21X1_388 ( .gnd(gnd), .vdd(vdd), .A(_5098_), .B(_4547__bF_buf54), .C(_5099_), .Y(_3673__9_) );
INVX1 INVX1_353 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__10_), .Y(_5100_) );
AOI22X1 AOI22X1_426 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[170]), .C(w_mem_inst_w_mem_10__10_), .D(_4548__bF_buf53), .Y(_5101_) );
OAI21X1 OAI21X1_389 ( .gnd(gnd), .vdd(vdd), .A(_5100_), .B(_4547__bF_buf53), .C(_5101_), .Y(_3673__10_) );
INVX1 INVX1_354 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__11_), .Y(_5102_) );
AOI22X1 AOI22X1_427 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[171]), .C(w_mem_inst_w_mem_10__11_), .D(_4548__bF_buf52), .Y(_5103_) );
OAI21X1 OAI21X1_390 ( .gnd(gnd), .vdd(vdd), .A(_5102_), .B(_4547__bF_buf52), .C(_5103_), .Y(_3673__11_) );
INVX1 INVX1_355 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__12_), .Y(_5104_) );
AOI22X1 AOI22X1_428 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[172]), .C(w_mem_inst_w_mem_10__12_), .D(_4548__bF_buf51), .Y(_5105_) );
OAI21X1 OAI21X1_391 ( .gnd(gnd), .vdd(vdd), .A(_5104_), .B(_4547__bF_buf51), .C(_5105_), .Y(_3673__12_) );
INVX1 INVX1_356 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__13_), .Y(_5106_) );
AOI22X1 AOI22X1_429 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[173]), .C(w_mem_inst_w_mem_10__13_), .D(_4548__bF_buf50), .Y(_5107_) );
OAI21X1 OAI21X1_392 ( .gnd(gnd), .vdd(vdd), .A(_5106_), .B(_4547__bF_buf50), .C(_5107_), .Y(_3673__13_) );
INVX1 INVX1_357 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__14_), .Y(_5108_) );
AOI22X1 AOI22X1_430 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[174]), .C(w_mem_inst_w_mem_10__14_), .D(_4548__bF_buf49), .Y(_5109_) );
OAI21X1 OAI21X1_393 ( .gnd(gnd), .vdd(vdd), .A(_5108_), .B(_4547__bF_buf49), .C(_5109_), .Y(_3673__14_) );
INVX1 INVX1_358 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__15_), .Y(_5110_) );
AOI22X1 AOI22X1_431 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[175]), .C(w_mem_inst_w_mem_10__15_), .D(_4548__bF_buf48), .Y(_5111_) );
OAI21X1 OAI21X1_394 ( .gnd(gnd), .vdd(vdd), .A(_5110_), .B(_4547__bF_buf48), .C(_5111_), .Y(_3673__15_) );
INVX1 INVX1_359 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__16_), .Y(_5112_) );
AOI22X1 AOI22X1_432 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[176]), .C(w_mem_inst_w_mem_10__16_), .D(_4548__bF_buf47), .Y(_5113_) );
OAI21X1 OAI21X1_395 ( .gnd(gnd), .vdd(vdd), .A(_5112_), .B(_4547__bF_buf47), .C(_5113_), .Y(_3673__16_) );
INVX1 INVX1_360 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__17_), .Y(_5114_) );
AOI22X1 AOI22X1_433 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[177]), .C(w_mem_inst_w_mem_10__17_), .D(_4548__bF_buf46), .Y(_5115_) );
OAI21X1 OAI21X1_396 ( .gnd(gnd), .vdd(vdd), .A(_5114_), .B(_4547__bF_buf46), .C(_5115_), .Y(_3673__17_) );
INVX1 INVX1_361 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__18_), .Y(_5116_) );
AOI22X1 AOI22X1_434 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[178]), .C(w_mem_inst_w_mem_10__18_), .D(_4548__bF_buf45), .Y(_5117_) );
OAI21X1 OAI21X1_397 ( .gnd(gnd), .vdd(vdd), .A(_5116_), .B(_4547__bF_buf45), .C(_5117_), .Y(_3673__18_) );
INVX1 INVX1_362 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__19_), .Y(_5118_) );
AOI22X1 AOI22X1_435 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[179]), .C(w_mem_inst_w_mem_10__19_), .D(_4548__bF_buf44), .Y(_5119_) );
OAI21X1 OAI21X1_398 ( .gnd(gnd), .vdd(vdd), .A(_5118_), .B(_4547__bF_buf44), .C(_5119_), .Y(_3673__19_) );
INVX1 INVX1_363 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__20_), .Y(_5120_) );
AOI22X1 AOI22X1_436 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[180]), .C(w_mem_inst_w_mem_10__20_), .D(_4548__bF_buf43), .Y(_5121_) );
OAI21X1 OAI21X1_399 ( .gnd(gnd), .vdd(vdd), .A(_5120_), .B(_4547__bF_buf43), .C(_5121_), .Y(_3673__20_) );
INVX1 INVX1_364 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__21_), .Y(_5122_) );
AOI22X1 AOI22X1_437 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[181]), .C(w_mem_inst_w_mem_10__21_), .D(_4548__bF_buf42), .Y(_5123_) );
OAI21X1 OAI21X1_400 ( .gnd(gnd), .vdd(vdd), .A(_5122_), .B(_4547__bF_buf42), .C(_5123_), .Y(_3673__21_) );
INVX1 INVX1_365 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__22_), .Y(_5124_) );
AOI22X1 AOI22X1_438 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[182]), .C(w_mem_inst_w_mem_10__22_), .D(_4548__bF_buf41), .Y(_5125_) );
OAI21X1 OAI21X1_401 ( .gnd(gnd), .vdd(vdd), .A(_5124_), .B(_4547__bF_buf41), .C(_5125_), .Y(_3673__22_) );
INVX1 INVX1_366 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__23_), .Y(_5126_) );
AOI22X1 AOI22X1_439 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[183]), .C(w_mem_inst_w_mem_10__23_), .D(_4548__bF_buf40), .Y(_5127_) );
OAI21X1 OAI21X1_402 ( .gnd(gnd), .vdd(vdd), .A(_5126_), .B(_4547__bF_buf40), .C(_5127_), .Y(_3673__23_) );
INVX1 INVX1_367 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__24_), .Y(_5128_) );
AOI22X1 AOI22X1_440 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[184]), .C(w_mem_inst_w_mem_10__24_), .D(_4548__bF_buf39), .Y(_5129_) );
OAI21X1 OAI21X1_403 ( .gnd(gnd), .vdd(vdd), .A(_5128_), .B(_4547__bF_buf39), .C(_5129_), .Y(_3673__24_) );
INVX1 INVX1_368 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__25_), .Y(_5130_) );
AOI22X1 AOI22X1_441 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[185]), .C(w_mem_inst_w_mem_10__25_), .D(_4548__bF_buf38), .Y(_5131_) );
OAI21X1 OAI21X1_404 ( .gnd(gnd), .vdd(vdd), .A(_5130_), .B(_4547__bF_buf38), .C(_5131_), .Y(_3673__25_) );
INVX1 INVX1_369 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__26_), .Y(_5132_) );
AOI22X1 AOI22X1_442 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[186]), .C(w_mem_inst_w_mem_10__26_), .D(_4548__bF_buf37), .Y(_5133_) );
OAI21X1 OAI21X1_405 ( .gnd(gnd), .vdd(vdd), .A(_5132_), .B(_4547__bF_buf37), .C(_5133_), .Y(_3673__26_) );
INVX1 INVX1_370 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__27_), .Y(_5134_) );
AOI22X1 AOI22X1_443 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[187]), .C(w_mem_inst_w_mem_10__27_), .D(_4548__bF_buf36), .Y(_5135_) );
OAI21X1 OAI21X1_406 ( .gnd(gnd), .vdd(vdd), .A(_5134_), .B(_4547__bF_buf36), .C(_5135_), .Y(_3673__27_) );
INVX1 INVX1_371 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__28_), .Y(_5136_) );
AOI22X1 AOI22X1_444 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[188]), .C(w_mem_inst_w_mem_10__28_), .D(_4548__bF_buf35), .Y(_5137_) );
OAI21X1 OAI21X1_407 ( .gnd(gnd), .vdd(vdd), .A(_5136_), .B(_4547__bF_buf35), .C(_5137_), .Y(_3673__28_) );
INVX1 INVX1_372 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__29_), .Y(_5138_) );
AOI22X1 AOI22X1_445 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[189]), .C(w_mem_inst_w_mem_10__29_), .D(_4548__bF_buf34), .Y(_5139_) );
OAI21X1 OAI21X1_408 ( .gnd(gnd), .vdd(vdd), .A(_5138_), .B(_4547__bF_buf34), .C(_5139_), .Y(_3673__29_) );
INVX1 INVX1_373 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__30_), .Y(_5140_) );
AOI22X1 AOI22X1_446 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[190]), .C(w_mem_inst_w_mem_10__30_), .D(_4548__bF_buf33), .Y(_5141_) );
OAI21X1 OAI21X1_409 ( .gnd(gnd), .vdd(vdd), .A(_5140_), .B(_4547__bF_buf33), .C(_5141_), .Y(_3673__30_) );
INVX1 INVX1_374 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__31_), .Y(_5142_) );
AOI22X1 AOI22X1_447 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[191]), .C(w_mem_inst_w_mem_10__31_), .D(_4548__bF_buf32), .Y(_5143_) );
OAI21X1 OAI21X1_410 ( .gnd(gnd), .vdd(vdd), .A(_5142_), .B(_4547__bF_buf32), .C(_5143_), .Y(_3673__31_) );
INVX1 INVX1_375 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__0_), .Y(_5144_) );
AOI22X1 AOI22X1_448 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[128]), .C(w_mem_inst_w_mem_11__0_), .D(_4548__bF_buf31), .Y(_5145_) );
OAI21X1 OAI21X1_411 ( .gnd(gnd), .vdd(vdd), .A(_5144_), .B(_4547__bF_buf31), .C(_5145_), .Y(_3674__0_) );
INVX1 INVX1_376 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__1_), .Y(_5146_) );
AOI22X1 AOI22X1_449 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[129]), .C(w_mem_inst_w_mem_11__1_), .D(_4548__bF_buf30), .Y(_5147_) );
OAI21X1 OAI21X1_412 ( .gnd(gnd), .vdd(vdd), .A(_5146_), .B(_4547__bF_buf30), .C(_5147_), .Y(_3674__1_) );
INVX1 INVX1_377 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__2_), .Y(_5148_) );
AOI22X1 AOI22X1_450 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[130]), .C(w_mem_inst_w_mem_11__2_), .D(_4548__bF_buf29), .Y(_5149_) );
OAI21X1 OAI21X1_413 ( .gnd(gnd), .vdd(vdd), .A(_5148_), .B(_4547__bF_buf29), .C(_5149_), .Y(_3674__2_) );
INVX1 INVX1_378 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__3_), .Y(_5150_) );
AOI22X1 AOI22X1_451 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[131]), .C(w_mem_inst_w_mem_11__3_), .D(_4548__bF_buf28), .Y(_5151_) );
OAI21X1 OAI21X1_414 ( .gnd(gnd), .vdd(vdd), .A(_5150_), .B(_4547__bF_buf28), .C(_5151_), .Y(_3674__3_) );
INVX1 INVX1_379 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__4_), .Y(_5152_) );
AOI22X1 AOI22X1_452 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[132]), .C(w_mem_inst_w_mem_11__4_), .D(_4548__bF_buf27), .Y(_5153_) );
OAI21X1 OAI21X1_415 ( .gnd(gnd), .vdd(vdd), .A(_5152_), .B(_4547__bF_buf27), .C(_5153_), .Y(_3674__4_) );
INVX1 INVX1_380 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__5_), .Y(_5154_) );
AOI22X1 AOI22X1_453 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[133]), .C(w_mem_inst_w_mem_11__5_), .D(_4548__bF_buf26), .Y(_5155_) );
OAI21X1 OAI21X1_416 ( .gnd(gnd), .vdd(vdd), .A(_5154_), .B(_4547__bF_buf26), .C(_5155_), .Y(_3674__5_) );
INVX1 INVX1_381 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__6_), .Y(_5156_) );
AOI22X1 AOI22X1_454 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[134]), .C(w_mem_inst_w_mem_11__6_), .D(_4548__bF_buf25), .Y(_5157_) );
OAI21X1 OAI21X1_417 ( .gnd(gnd), .vdd(vdd), .A(_5156_), .B(_4547__bF_buf25), .C(_5157_), .Y(_3674__6_) );
INVX1 INVX1_382 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__7_), .Y(_5158_) );
AOI22X1 AOI22X1_455 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[135]), .C(w_mem_inst_w_mem_11__7_), .D(_4548__bF_buf24), .Y(_5159_) );
OAI21X1 OAI21X1_418 ( .gnd(gnd), .vdd(vdd), .A(_5158_), .B(_4547__bF_buf24), .C(_5159_), .Y(_3674__7_) );
INVX1 INVX1_383 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__8_), .Y(_5160_) );
AOI22X1 AOI22X1_456 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[136]), .C(w_mem_inst_w_mem_11__8_), .D(_4548__bF_buf23), .Y(_5161_) );
OAI21X1 OAI21X1_419 ( .gnd(gnd), .vdd(vdd), .A(_5160_), .B(_4547__bF_buf23), .C(_5161_), .Y(_3674__8_) );
INVX1 INVX1_384 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__9_), .Y(_5162_) );
AOI22X1 AOI22X1_457 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[137]), .C(w_mem_inst_w_mem_11__9_), .D(_4548__bF_buf22), .Y(_5163_) );
OAI21X1 OAI21X1_420 ( .gnd(gnd), .vdd(vdd), .A(_5162_), .B(_4547__bF_buf22), .C(_5163_), .Y(_3674__9_) );
INVX1 INVX1_385 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__10_), .Y(_5164_) );
AOI22X1 AOI22X1_458 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[138]), .C(w_mem_inst_w_mem_11__10_), .D(_4548__bF_buf21), .Y(_5165_) );
OAI21X1 OAI21X1_421 ( .gnd(gnd), .vdd(vdd), .A(_5164_), .B(_4547__bF_buf21), .C(_5165_), .Y(_3674__10_) );
INVX1 INVX1_386 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__11_), .Y(_5166_) );
AOI22X1 AOI22X1_459 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[139]), .C(w_mem_inst_w_mem_11__11_), .D(_4548__bF_buf20), .Y(_5167_) );
OAI21X1 OAI21X1_422 ( .gnd(gnd), .vdd(vdd), .A(_5166_), .B(_4547__bF_buf20), .C(_5167_), .Y(_3674__11_) );
INVX1 INVX1_387 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__12_), .Y(_5168_) );
AOI22X1 AOI22X1_460 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[140]), .C(w_mem_inst_w_mem_11__12_), .D(_4548__bF_buf19), .Y(_5169_) );
OAI21X1 OAI21X1_423 ( .gnd(gnd), .vdd(vdd), .A(_5168_), .B(_4547__bF_buf19), .C(_5169_), .Y(_3674__12_) );
INVX1 INVX1_388 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__13_), .Y(_5170_) );
AOI22X1 AOI22X1_461 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[141]), .C(w_mem_inst_w_mem_11__13_), .D(_4548__bF_buf18), .Y(_5171_) );
OAI21X1 OAI21X1_424 ( .gnd(gnd), .vdd(vdd), .A(_5170_), .B(_4547__bF_buf18), .C(_5171_), .Y(_3674__13_) );
INVX1 INVX1_389 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__14_), .Y(_5172_) );
AOI22X1 AOI22X1_462 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[142]), .C(w_mem_inst_w_mem_11__14_), .D(_4548__bF_buf17), .Y(_5173_) );
OAI21X1 OAI21X1_425 ( .gnd(gnd), .vdd(vdd), .A(_5172_), .B(_4547__bF_buf17), .C(_5173_), .Y(_3674__14_) );
INVX1 INVX1_390 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__15_), .Y(_5174_) );
AOI22X1 AOI22X1_463 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[143]), .C(w_mem_inst_w_mem_11__15_), .D(_4548__bF_buf16), .Y(_5175_) );
OAI21X1 OAI21X1_426 ( .gnd(gnd), .vdd(vdd), .A(_5174_), .B(_4547__bF_buf16), .C(_5175_), .Y(_3674__15_) );
INVX1 INVX1_391 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__16_), .Y(_5176_) );
AOI22X1 AOI22X1_464 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[144]), .C(w_mem_inst_w_mem_11__16_), .D(_4548__bF_buf15), .Y(_5177_) );
OAI21X1 OAI21X1_427 ( .gnd(gnd), .vdd(vdd), .A(_5176_), .B(_4547__bF_buf15), .C(_5177_), .Y(_3674__16_) );
INVX1 INVX1_392 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__17_), .Y(_5178_) );
AOI22X1 AOI22X1_465 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[145]), .C(w_mem_inst_w_mem_11__17_), .D(_4548__bF_buf14), .Y(_5179_) );
OAI21X1 OAI21X1_428 ( .gnd(gnd), .vdd(vdd), .A(_5178_), .B(_4547__bF_buf14), .C(_5179_), .Y(_3674__17_) );
INVX1 INVX1_393 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__18_), .Y(_5180_) );
AOI22X1 AOI22X1_466 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[146]), .C(w_mem_inst_w_mem_11__18_), .D(_4548__bF_buf13), .Y(_5181_) );
OAI21X1 OAI21X1_429 ( .gnd(gnd), .vdd(vdd), .A(_5180_), .B(_4547__bF_buf13), .C(_5181_), .Y(_3674__18_) );
INVX1 INVX1_394 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__19_), .Y(_5182_) );
AOI22X1 AOI22X1_467 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[147]), .C(w_mem_inst_w_mem_11__19_), .D(_4548__bF_buf12), .Y(_5183_) );
OAI21X1 OAI21X1_430 ( .gnd(gnd), .vdd(vdd), .A(_5182_), .B(_4547__bF_buf12), .C(_5183_), .Y(_3674__19_) );
INVX1 INVX1_395 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__20_), .Y(_5184_) );
AOI22X1 AOI22X1_468 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[148]), .C(w_mem_inst_w_mem_11__20_), .D(_4548__bF_buf11), .Y(_5185_) );
OAI21X1 OAI21X1_431 ( .gnd(gnd), .vdd(vdd), .A(_5184_), .B(_4547__bF_buf11), .C(_5185_), .Y(_3674__20_) );
INVX1 INVX1_396 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__21_), .Y(_5186_) );
AOI22X1 AOI22X1_469 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[149]), .C(w_mem_inst_w_mem_11__21_), .D(_4548__bF_buf10), .Y(_5187_) );
OAI21X1 OAI21X1_432 ( .gnd(gnd), .vdd(vdd), .A(_5186_), .B(_4547__bF_buf10), .C(_5187_), .Y(_3674__21_) );
INVX1 INVX1_397 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__22_), .Y(_5188_) );
AOI22X1 AOI22X1_470 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[150]), .C(w_mem_inst_w_mem_11__22_), .D(_4548__bF_buf9), .Y(_5189_) );
OAI21X1 OAI21X1_433 ( .gnd(gnd), .vdd(vdd), .A(_5188_), .B(_4547__bF_buf9), .C(_5189_), .Y(_3674__22_) );
INVX1 INVX1_398 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__23_), .Y(_5190_) );
AOI22X1 AOI22X1_471 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[151]), .C(w_mem_inst_w_mem_11__23_), .D(_4548__bF_buf8), .Y(_5191_) );
OAI21X1 OAI21X1_434 ( .gnd(gnd), .vdd(vdd), .A(_5190_), .B(_4547__bF_buf8), .C(_5191_), .Y(_3674__23_) );
INVX1 INVX1_399 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__24_), .Y(_5192_) );
AOI22X1 AOI22X1_472 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[152]), .C(w_mem_inst_w_mem_11__24_), .D(_4548__bF_buf7), .Y(_5193_) );
OAI21X1 OAI21X1_435 ( .gnd(gnd), .vdd(vdd), .A(_5192_), .B(_4547__bF_buf7), .C(_5193_), .Y(_3674__24_) );
INVX1 INVX1_400 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__25_), .Y(_5194_) );
AOI22X1 AOI22X1_473 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[153]), .C(w_mem_inst_w_mem_11__25_), .D(_4548__bF_buf6), .Y(_5195_) );
OAI21X1 OAI21X1_436 ( .gnd(gnd), .vdd(vdd), .A(_5194_), .B(_4547__bF_buf6), .C(_5195_), .Y(_3674__25_) );
INVX1 INVX1_401 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__26_), .Y(_5196_) );
AOI22X1 AOI22X1_474 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[154]), .C(w_mem_inst_w_mem_11__26_), .D(_4548__bF_buf5), .Y(_5197_) );
OAI21X1 OAI21X1_437 ( .gnd(gnd), .vdd(vdd), .A(_5196_), .B(_4547__bF_buf5), .C(_5197_), .Y(_3674__26_) );
INVX1 INVX1_402 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__27_), .Y(_5198_) );
AOI22X1 AOI22X1_475 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[155]), .C(w_mem_inst_w_mem_11__27_), .D(_4548__bF_buf4), .Y(_5199_) );
OAI21X1 OAI21X1_438 ( .gnd(gnd), .vdd(vdd), .A(_5198_), .B(_4547__bF_buf4), .C(_5199_), .Y(_3674__27_) );
INVX1 INVX1_403 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__28_), .Y(_5200_) );
AOI22X1 AOI22X1_476 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[156]), .C(w_mem_inst_w_mem_11__28_), .D(_4548__bF_buf3), .Y(_5201_) );
OAI21X1 OAI21X1_439 ( .gnd(gnd), .vdd(vdd), .A(_5200_), .B(_4547__bF_buf3), .C(_5201_), .Y(_3674__28_) );
INVX1 INVX1_404 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__29_), .Y(_5202_) );
AOI22X1 AOI22X1_477 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[157]), .C(w_mem_inst_w_mem_11__29_), .D(_4548__bF_buf2), .Y(_5203_) );
OAI21X1 OAI21X1_440 ( .gnd(gnd), .vdd(vdd), .A(_5202_), .B(_4547__bF_buf2), .C(_5203_), .Y(_3674__29_) );
INVX1 INVX1_405 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__30_), .Y(_5204_) );
AOI22X1 AOI22X1_478 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[158]), .C(w_mem_inst_w_mem_11__30_), .D(_4548__bF_buf1), .Y(_5205_) );
OAI21X1 OAI21X1_441 ( .gnd(gnd), .vdd(vdd), .A(_5204_), .B(_4547__bF_buf1), .C(_5205_), .Y(_3674__30_) );
INVX1 INVX1_406 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__31_), .Y(_5206_) );
AOI22X1 AOI22X1_479 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[159]), .C(w_mem_inst_w_mem_11__31_), .D(_4548__bF_buf0), .Y(_5207_) );
OAI21X1 OAI21X1_442 ( .gnd(gnd), .vdd(vdd), .A(_5206_), .B(_4547__bF_buf0), .C(_5207_), .Y(_3674__31_) );
AOI22X1 AOI22X1_480 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[96]), .C(w_mem_inst_w_mem_12__0_), .D(_4548__bF_buf63), .Y(_5208_) );
OAI21X1 OAI21X1_443 ( .gnd(gnd), .vdd(vdd), .A(_3714_), .B(_4547__bF_buf63), .C(_5208_), .Y(_3675__0_) );
AOI22X1 AOI22X1_481 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[97]), .C(w_mem_inst_w_mem_12__1_), .D(_4548__bF_buf62), .Y(_5209_) );
OAI21X1 OAI21X1_444 ( .gnd(gnd), .vdd(vdd), .A(_3758_), .B(_4547__bF_buf62), .C(_5209_), .Y(_3675__1_) );
INVX1 INVX1_407 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__2_), .Y(_5210_) );
AOI22X1 AOI22X1_482 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[98]), .C(w_mem_inst_w_mem_12__2_), .D(_4548__bF_buf61), .Y(_5211_) );
OAI21X1 OAI21X1_445 ( .gnd(gnd), .vdd(vdd), .A(_5210_), .B(_4547__bF_buf61), .C(_5211_), .Y(_3675__2_) );
AOI22X1 AOI22X1_483 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[99]), .C(w_mem_inst_w_mem_12__3_), .D(_4548__bF_buf60), .Y(_5212_) );
OAI21X1 OAI21X1_446 ( .gnd(gnd), .vdd(vdd), .A(_3810_), .B(_4547__bF_buf60), .C(_5212_), .Y(_3675__3_) );
INVX1 INVX1_408 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__4_), .Y(_5213_) );
AOI22X1 AOI22X1_484 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[100]), .C(w_mem_inst_w_mem_12__4_), .D(_4548__bF_buf59), .Y(_5214_) );
OAI21X1 OAI21X1_447 ( .gnd(gnd), .vdd(vdd), .A(_5213_), .B(_4547__bF_buf59), .C(_5214_), .Y(_3675__4_) );
INVX1 INVX1_409 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__5_), .Y(_5215_) );
AOI22X1 AOI22X1_485 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[101]), .C(w_mem_inst_w_mem_12__5_), .D(_4548__bF_buf58), .Y(_5216_) );
OAI21X1 OAI21X1_448 ( .gnd(gnd), .vdd(vdd), .A(_5215_), .B(_4547__bF_buf58), .C(_5216_), .Y(_3675__5_) );
AOI22X1 AOI22X1_486 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[102]), .C(w_mem_inst_w_mem_12__6_), .D(_4548__bF_buf57), .Y(_5217_) );
OAI21X1 OAI21X1_449 ( .gnd(gnd), .vdd(vdd), .A(_3890_), .B(_4547__bF_buf57), .C(_5217_), .Y(_3675__6_) );
AOI22X1 AOI22X1_487 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[103]), .C(w_mem_inst_w_mem_12__7_), .D(_4548__bF_buf56), .Y(_5218_) );
OAI21X1 OAI21X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3911_), .B(_4547__bF_buf56), .C(_5218_), .Y(_3675__7_) );
INVX1 INVX1_410 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__8_), .Y(_5219_) );
AOI22X1 AOI22X1_488 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[104]), .C(w_mem_inst_w_mem_12__8_), .D(_4548__bF_buf55), .Y(_5220_) );
OAI21X1 OAI21X1_451 ( .gnd(gnd), .vdd(vdd), .A(_5219_), .B(_4547__bF_buf55), .C(_5220_), .Y(_3675__8_) );
AOI22X1 AOI22X1_489 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[105]), .C(w_mem_inst_w_mem_12__9_), .D(_4548__bF_buf54), .Y(_5221_) );
OAI21X1 OAI21X1_452 ( .gnd(gnd), .vdd(vdd), .A(_3964_), .B(_4547__bF_buf54), .C(_5221_), .Y(_3675__9_) );
AOI22X1 AOI22X1_490 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[106]), .C(w_mem_inst_w_mem_12__10_), .D(_4548__bF_buf53), .Y(_5222_) );
OAI21X1 OAI21X1_453 ( .gnd(gnd), .vdd(vdd), .A(_3989_), .B(_4547__bF_buf53), .C(_5222_), .Y(_3675__10_) );
AOI22X1 AOI22X1_491 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[107]), .C(w_mem_inst_w_mem_12__11_), .D(_4548__bF_buf52), .Y(_5223_) );
OAI21X1 OAI21X1_454 ( .gnd(gnd), .vdd(vdd), .A(_4014_), .B(_4547__bF_buf52), .C(_5223_), .Y(_3675__11_) );
AOI22X1 AOI22X1_492 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[108]), .C(w_mem_inst_w_mem_12__12_), .D(_4548__bF_buf51), .Y(_5224_) );
OAI21X1 OAI21X1_455 ( .gnd(gnd), .vdd(vdd), .A(_4038_), .B(_4547__bF_buf51), .C(_5224_), .Y(_3675__12_) );
AOI22X1 AOI22X1_493 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[109]), .C(w_mem_inst_w_mem_12__13_), .D(_4548__bF_buf50), .Y(_5225_) );
OAI21X1 OAI21X1_456 ( .gnd(gnd), .vdd(vdd), .A(_4064_), .B(_4547__bF_buf50), .C(_5225_), .Y(_3675__13_) );
AOI22X1 AOI22X1_494 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[110]), .C(w_mem_inst_w_mem_12__14_), .D(_4548__bF_buf49), .Y(_5226_) );
OAI21X1 OAI21X1_457 ( .gnd(gnd), .vdd(vdd), .A(_4088_), .B(_4547__bF_buf49), .C(_5226_), .Y(_3675__14_) );
AOI22X1 AOI22X1_495 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[111]), .C(w_mem_inst_w_mem_12__15_), .D(_4548__bF_buf48), .Y(_5227_) );
OAI21X1 OAI21X1_458 ( .gnd(gnd), .vdd(vdd), .A(_4109_), .B(_4547__bF_buf48), .C(_5227_), .Y(_3675__15_) );
INVX1 INVX1_411 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__16_), .Y(_5228_) );
AOI22X1 AOI22X1_496 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[112]), .C(w_mem_inst_w_mem_12__16_), .D(_4548__bF_buf47), .Y(_5229_) );
OAI21X1 OAI21X1_459 ( .gnd(gnd), .vdd(vdd), .A(_5228_), .B(_4547__bF_buf47), .C(_5229_), .Y(_3675__16_) );
AOI22X1 AOI22X1_497 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[113]), .C(w_mem_inst_w_mem_12__17_), .D(_4548__bF_buf46), .Y(_5230_) );
OAI21X1 OAI21X1_460 ( .gnd(gnd), .vdd(vdd), .A(_4162_), .B(_4547__bF_buf46), .C(_5230_), .Y(_3675__17_) );
AOI22X1 AOI22X1_498 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[114]), .C(w_mem_inst_w_mem_12__18_), .D(_4548__bF_buf45), .Y(_5231_) );
OAI21X1 OAI21X1_461 ( .gnd(gnd), .vdd(vdd), .A(_4187_), .B(_4547__bF_buf45), .C(_5231_), .Y(_3675__18_) );
AOI22X1 AOI22X1_499 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[115]), .C(w_mem_inst_w_mem_12__19_), .D(_4548__bF_buf44), .Y(_5232_) );
OAI21X1 OAI21X1_462 ( .gnd(gnd), .vdd(vdd), .A(_4212_), .B(_4547__bF_buf44), .C(_5232_), .Y(_3675__19_) );
AOI22X1 AOI22X1_500 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[116]), .C(w_mem_inst_w_mem_12__20_), .D(_4548__bF_buf43), .Y(_5233_) );
OAI21X1 OAI21X1_463 ( .gnd(gnd), .vdd(vdd), .A(_4236_), .B(_4547__bF_buf43), .C(_5233_), .Y(_3675__20_) );
AOI22X1 AOI22X1_501 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[117]), .C(w_mem_inst_w_mem_12__21_), .D(_4548__bF_buf42), .Y(_5234_) );
OAI21X1 OAI21X1_464 ( .gnd(gnd), .vdd(vdd), .A(_4262_), .B(_4547__bF_buf42), .C(_5234_), .Y(_3675__21_) );
AOI22X1 AOI22X1_502 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[118]), .C(w_mem_inst_w_mem_12__22_), .D(_4548__bF_buf41), .Y(_5235_) );
OAI21X1 OAI21X1_465 ( .gnd(gnd), .vdd(vdd), .A(_4286_), .B(_4547__bF_buf41), .C(_5235_), .Y(_3675__22_) );
AOI22X1 AOI22X1_503 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[119]), .C(w_mem_inst_w_mem_12__23_), .D(_4548__bF_buf40), .Y(_5236_) );
OAI21X1 OAI21X1_466 ( .gnd(gnd), .vdd(vdd), .A(_4307_), .B(_4547__bF_buf40), .C(_5236_), .Y(_3675__23_) );
INVX1 INVX1_412 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__24_), .Y(_5237_) );
AOI22X1 AOI22X1_504 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[120]), .C(w_mem_inst_w_mem_12__24_), .D(_4548__bF_buf39), .Y(_5238_) );
OAI21X1 OAI21X1_467 ( .gnd(gnd), .vdd(vdd), .A(_5237_), .B(_4547__bF_buf39), .C(_5238_), .Y(_3675__24_) );
AOI22X1 AOI22X1_505 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[121]), .C(w_mem_inst_w_mem_12__25_), .D(_4548__bF_buf38), .Y(_5239_) );
OAI21X1 OAI21X1_468 ( .gnd(gnd), .vdd(vdd), .A(_4360_), .B(_4547__bF_buf38), .C(_5239_), .Y(_3675__25_) );
AOI22X1 AOI22X1_506 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[122]), .C(w_mem_inst_w_mem_12__26_), .D(_4548__bF_buf37), .Y(_5240_) );
OAI21X1 OAI21X1_469 ( .gnd(gnd), .vdd(vdd), .A(_4385_), .B(_4547__bF_buf37), .C(_5240_), .Y(_3675__26_) );
AOI22X1 AOI22X1_507 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[123]), .C(w_mem_inst_w_mem_12__27_), .D(_4548__bF_buf36), .Y(_5241_) );
OAI21X1 OAI21X1_470 ( .gnd(gnd), .vdd(vdd), .A(_4410_), .B(_4547__bF_buf36), .C(_5241_), .Y(_3675__27_) );
AOI22X1 AOI22X1_508 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[124]), .C(w_mem_inst_w_mem_12__28_), .D(_4548__bF_buf35), .Y(_5242_) );
OAI21X1 OAI21X1_471 ( .gnd(gnd), .vdd(vdd), .A(_4434_), .B(_4547__bF_buf35), .C(_5242_), .Y(_3675__28_) );
AOI22X1 AOI22X1_509 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[125]), .C(w_mem_inst_w_mem_12__29_), .D(_4548__bF_buf34), .Y(_5243_) );
OAI21X1 OAI21X1_472 ( .gnd(gnd), .vdd(vdd), .A(_4460_), .B(_4547__bF_buf34), .C(_5243_), .Y(_3675__29_) );
AOI22X1 AOI22X1_510 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[126]), .C(w_mem_inst_w_mem_12__30_), .D(_4548__bF_buf33), .Y(_5244_) );
OAI21X1 OAI21X1_473 ( .gnd(gnd), .vdd(vdd), .A(_4484_), .B(_4547__bF_buf33), .C(_5244_), .Y(_3675__30_) );
INVX1 INVX1_413 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__31_), .Y(_5245_) );
AOI22X1 AOI22X1_511 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[127]), .C(w_mem_inst_w_mem_12__31_), .D(_4548__bF_buf32), .Y(_5246_) );
OAI21X1 OAI21X1_474 ( .gnd(gnd), .vdd(vdd), .A(_5245_), .B(_4547__bF_buf32), .C(_5246_), .Y(_3675__31_) );
INVX1 INVX1_414 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__0_), .Y(_5247_) );
AOI22X1 AOI22X1_512 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[64]), .C(w_mem_inst_w_mem_13__0_), .D(_4548__bF_buf31), .Y(_5248_) );
OAI21X1 OAI21X1_475 ( .gnd(gnd), .vdd(vdd), .A(_5247_), .B(_4547__bF_buf31), .C(_5248_), .Y(_3676__0_) );
INVX1 INVX1_415 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__1_), .Y(_5249_) );
AOI22X1 AOI22X1_513 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[65]), .C(w_mem_inst_w_mem_13__1_), .D(_4548__bF_buf30), .Y(_5250_) );
OAI21X1 OAI21X1_476 ( .gnd(gnd), .vdd(vdd), .A(_5249_), .B(_4547__bF_buf30), .C(_5250_), .Y(_3676__1_) );
INVX1 INVX1_416 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__2_), .Y(_5251_) );
AOI22X1 AOI22X1_514 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[66]), .C(w_mem_inst_w_mem_13__2_), .D(_4548__bF_buf29), .Y(_5252_) );
OAI21X1 OAI21X1_477 ( .gnd(gnd), .vdd(vdd), .A(_5251_), .B(_4547__bF_buf29), .C(_5252_), .Y(_3676__2_) );
INVX1 INVX1_417 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__3_), .Y(_5253_) );
AOI22X1 AOI22X1_515 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[67]), .C(w_mem_inst_w_mem_13__3_), .D(_4548__bF_buf28), .Y(_5254_) );
OAI21X1 OAI21X1_478 ( .gnd(gnd), .vdd(vdd), .A(_5253_), .B(_4547__bF_buf28), .C(_5254_), .Y(_3676__3_) );
AOI22X1 AOI22X1_516 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[68]), .C(w_mem_inst_w_mem_13__4_), .D(_4548__bF_buf27), .Y(_5255_) );
OAI21X1 OAI21X1_479 ( .gnd(gnd), .vdd(vdd), .A(_3836_), .B(_4547__bF_buf27), .C(_5255_), .Y(_3676__4_) );
INVX1 INVX1_418 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__5_), .Y(_5256_) );
AOI22X1 AOI22X1_517 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[69]), .C(w_mem_inst_w_mem_13__5_), .D(_4548__bF_buf26), .Y(_5257_) );
OAI21X1 OAI21X1_480 ( .gnd(gnd), .vdd(vdd), .A(_5256_), .B(_4547__bF_buf26), .C(_5257_), .Y(_3676__5_) );
AOI22X1 AOI22X1_518 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[70]), .C(w_mem_inst_w_mem_13__6_), .D(_4548__bF_buf25), .Y(_5258_) );
OAI21X1 OAI21X1_481 ( .gnd(gnd), .vdd(vdd), .A(_3885_), .B(_4547__bF_buf25), .C(_5258_), .Y(_3676__6_) );
INVX1 INVX1_419 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__7_), .Y(_5259_) );
AOI22X1 AOI22X1_519 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[71]), .C(w_mem_inst_w_mem_13__7_), .D(_4548__bF_buf24), .Y(_5260_) );
OAI21X1 OAI21X1_482 ( .gnd(gnd), .vdd(vdd), .A(_5259_), .B(_4547__bF_buf24), .C(_5260_), .Y(_3676__7_) );
INVX1 INVX1_420 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__8_), .Y(_5261_) );
AOI22X1 AOI22X1_520 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[72]), .C(w_mem_inst_w_mem_13__8_), .D(_4548__bF_buf23), .Y(_5262_) );
OAI21X1 OAI21X1_483 ( .gnd(gnd), .vdd(vdd), .A(_5261_), .B(_4547__bF_buf23), .C(_5262_), .Y(_3676__8_) );
INVX1 INVX1_421 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__9_), .Y(_5263_) );
AOI22X1 AOI22X1_521 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[73]), .C(w_mem_inst_w_mem_13__9_), .D(_4548__bF_buf22), .Y(_5264_) );
OAI21X1 OAI21X1_484 ( .gnd(gnd), .vdd(vdd), .A(_5263_), .B(_4547__bF_buf22), .C(_5264_), .Y(_3676__9_) );
INVX1 INVX1_422 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__10_), .Y(_5265_) );
AOI22X1 AOI22X1_522 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[74]), .C(w_mem_inst_w_mem_13__10_), .D(_4548__bF_buf21), .Y(_5266_) );
OAI21X1 OAI21X1_485 ( .gnd(gnd), .vdd(vdd), .A(_5265_), .B(_4547__bF_buf21), .C(_5266_), .Y(_3676__10_) );
INVX1 INVX1_423 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__11_), .Y(_5267_) );
AOI22X1 AOI22X1_523 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[75]), .C(w_mem_inst_w_mem_13__11_), .D(_4548__bF_buf20), .Y(_5268_) );
OAI21X1 OAI21X1_486 ( .gnd(gnd), .vdd(vdd), .A(_5267_), .B(_4547__bF_buf20), .C(_5268_), .Y(_3676__11_) );
INVX1 INVX1_424 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__12_), .Y(_5269_) );
AOI22X1 AOI22X1_524 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[76]), .C(w_mem_inst_w_mem_13__12_), .D(_4548__bF_buf19), .Y(_5270_) );
OAI21X1 OAI21X1_487 ( .gnd(gnd), .vdd(vdd), .A(_5269_), .B(_4547__bF_buf19), .C(_5270_), .Y(_3676__12_) );
INVX1 INVX1_425 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__13_), .Y(_5271_) );
AOI22X1 AOI22X1_525 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[77]), .C(w_mem_inst_w_mem_13__13_), .D(_4548__bF_buf18), .Y(_5272_) );
OAI21X1 OAI21X1_488 ( .gnd(gnd), .vdd(vdd), .A(_5271_), .B(_4547__bF_buf18), .C(_5272_), .Y(_3676__13_) );
AOI22X1 AOI22X1_526 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[78]), .C(w_mem_inst_w_mem_13__14_), .D(_4548__bF_buf17), .Y(_5273_) );
OAI21X1 OAI21X1_489 ( .gnd(gnd), .vdd(vdd), .A(_4083_), .B(_4547__bF_buf17), .C(_5273_), .Y(_3676__14_) );
INVX1 INVX1_426 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__15_), .Y(_5274_) );
AOI22X1 AOI22X1_527 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[79]), .C(w_mem_inst_w_mem_13__15_), .D(_4548__bF_buf16), .Y(_5275_) );
OAI21X1 OAI21X1_490 ( .gnd(gnd), .vdd(vdd), .A(_5274_), .B(_4547__bF_buf16), .C(_5275_), .Y(_3676__15_) );
INVX1 INVX1_427 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__16_), .Y(_5276_) );
AOI22X1 AOI22X1_528 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[80]), .C(w_mem_inst_w_mem_13__16_), .D(_4548__bF_buf15), .Y(_5277_) );
OAI21X1 OAI21X1_491 ( .gnd(gnd), .vdd(vdd), .A(_5276_), .B(_4547__bF_buf15), .C(_5277_), .Y(_3676__16_) );
INVX1 INVX1_428 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__17_), .Y(_5278_) );
AOI22X1 AOI22X1_529 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[81]), .C(w_mem_inst_w_mem_13__17_), .D(_4548__bF_buf14), .Y(_5279_) );
OAI21X1 OAI21X1_492 ( .gnd(gnd), .vdd(vdd), .A(_5278_), .B(_4547__bF_buf14), .C(_5279_), .Y(_3676__17_) );
INVX1 INVX1_429 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__18_), .Y(_5280_) );
AOI22X1 AOI22X1_530 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[82]), .C(w_mem_inst_w_mem_13__18_), .D(_4548__bF_buf13), .Y(_5281_) );
OAI21X1 OAI21X1_493 ( .gnd(gnd), .vdd(vdd), .A(_5280_), .B(_4547__bF_buf13), .C(_5281_), .Y(_3676__18_) );
INVX1 INVX1_430 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__19_), .Y(_5282_) );
AOI22X1 AOI22X1_531 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[83]), .C(w_mem_inst_w_mem_13__19_), .D(_4548__bF_buf12), .Y(_5283_) );
OAI21X1 OAI21X1_494 ( .gnd(gnd), .vdd(vdd), .A(_5282_), .B(_4547__bF_buf12), .C(_5283_), .Y(_3676__19_) );
INVX1 INVX1_431 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__20_), .Y(_5284_) );
AOI22X1 AOI22X1_532 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[84]), .C(w_mem_inst_w_mem_13__20_), .D(_4548__bF_buf11), .Y(_5285_) );
OAI21X1 OAI21X1_495 ( .gnd(gnd), .vdd(vdd), .A(_5284_), .B(_4547__bF_buf11), .C(_5285_), .Y(_3676__20_) );
INVX1 INVX1_432 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__21_), .Y(_5286_) );
AOI22X1 AOI22X1_533 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[85]), .C(w_mem_inst_w_mem_13__21_), .D(_4548__bF_buf10), .Y(_5287_) );
OAI21X1 OAI21X1_496 ( .gnd(gnd), .vdd(vdd), .A(_5286_), .B(_4547__bF_buf10), .C(_5287_), .Y(_3676__21_) );
AOI22X1 AOI22X1_534 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[86]), .C(w_mem_inst_w_mem_13__22_), .D(_4548__bF_buf9), .Y(_5288_) );
OAI21X1 OAI21X1_497 ( .gnd(gnd), .vdd(vdd), .A(_4281_), .B(_4547__bF_buf9), .C(_5288_), .Y(_3676__22_) );
INVX1 INVX1_433 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__23_), .Y(_5289_) );
AOI22X1 AOI22X1_535 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[87]), .C(w_mem_inst_w_mem_13__23_), .D(_4548__bF_buf8), .Y(_5290_) );
OAI21X1 OAI21X1_498 ( .gnd(gnd), .vdd(vdd), .A(_5289_), .B(_4547__bF_buf8), .C(_5290_), .Y(_3676__23_) );
INVX1 INVX1_434 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__24_), .Y(_5291_) );
AOI22X1 AOI22X1_536 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[88]), .C(w_mem_inst_w_mem_13__24_), .D(_4548__bF_buf7), .Y(_5292_) );
OAI21X1 OAI21X1_499 ( .gnd(gnd), .vdd(vdd), .A(_5291_), .B(_4547__bF_buf7), .C(_5292_), .Y(_3676__24_) );
INVX1 INVX1_435 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__25_), .Y(_5293_) );
AOI22X1 AOI22X1_537 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[89]), .C(w_mem_inst_w_mem_13__25_), .D(_4548__bF_buf6), .Y(_5294_) );
OAI21X1 OAI21X1_500 ( .gnd(gnd), .vdd(vdd), .A(_5293_), .B(_4547__bF_buf6), .C(_5294_), .Y(_3676__25_) );
INVX1 INVX1_436 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__26_), .Y(_5295_) );
AOI22X1 AOI22X1_538 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[90]), .C(w_mem_inst_w_mem_13__26_), .D(_4548__bF_buf5), .Y(_5296_) );
OAI21X1 OAI21X1_501 ( .gnd(gnd), .vdd(vdd), .A(_5295_), .B(_4547__bF_buf5), .C(_5296_), .Y(_3676__26_) );
INVX1 INVX1_437 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__27_), .Y(_5297_) );
AOI22X1 AOI22X1_539 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[91]), .C(w_mem_inst_w_mem_13__27_), .D(_4548__bF_buf4), .Y(_5298_) );
OAI21X1 OAI21X1_502 ( .gnd(gnd), .vdd(vdd), .A(_5297_), .B(_4547__bF_buf4), .C(_5298_), .Y(_3676__27_) );
INVX1 INVX1_438 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__28_), .Y(_5299_) );
AOI22X1 AOI22X1_540 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[92]), .C(w_mem_inst_w_mem_13__28_), .D(_4548__bF_buf3), .Y(_5300_) );
OAI21X1 OAI21X1_503 ( .gnd(gnd), .vdd(vdd), .A(_5299_), .B(_4547__bF_buf3), .C(_5300_), .Y(_3676__28_) );
INVX1 INVX1_439 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__29_), .Y(_5301_) );
AOI22X1 AOI22X1_541 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[93]), .C(w_mem_inst_w_mem_13__29_), .D(_4548__bF_buf2), .Y(_5302_) );
OAI21X1 OAI21X1_504 ( .gnd(gnd), .vdd(vdd), .A(_5301_), .B(_4547__bF_buf2), .C(_5302_), .Y(_3676__29_) );
AOI22X1 AOI22X1_542 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[94]), .C(w_mem_inst_w_mem_13__30_), .D(_4548__bF_buf1), .Y(_5303_) );
OAI21X1 OAI21X1_505 ( .gnd(gnd), .vdd(vdd), .A(_4479_), .B(_4547__bF_buf1), .C(_5303_), .Y(_3676__30_) );
AOI22X1 AOI22X1_543 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[95]), .C(w_mem_inst_w_mem_13__31_), .D(_4548__bF_buf0), .Y(_5304_) );
OAI21X1 OAI21X1_506 ( .gnd(gnd), .vdd(vdd), .A(_4506_), .B(_4547__bF_buf0), .C(_5304_), .Y(_3676__31_) );
INVX1 INVX1_440 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__0_), .Y(_5305_) );
AOI22X1 AOI22X1_544 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf61), .B(block[32]), .C(w_mem_inst_w_mem_14__0_), .D(_4548__bF_buf63), .Y(_5306_) );
OAI21X1 OAI21X1_507 ( .gnd(gnd), .vdd(vdd), .A(_5305_), .B(_4547__bF_buf63), .C(_5306_), .Y(_3677__0_) );
INVX1 INVX1_441 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__1_), .Y(_5307_) );
AOI22X1 AOI22X1_545 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf60), .B(block[33]), .C(w_mem_inst_w_mem_14__1_), .D(_4548__bF_buf62), .Y(_5308_) );
OAI21X1 OAI21X1_508 ( .gnd(gnd), .vdd(vdd), .A(_5307_), .B(_4547__bF_buf62), .C(_5308_), .Y(_3677__1_) );
INVX1 INVX1_442 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__2_), .Y(_5309_) );
AOI22X1 AOI22X1_546 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf59), .B(block[34]), .C(w_mem_inst_w_mem_14__2_), .D(_4548__bF_buf61), .Y(_5310_) );
OAI21X1 OAI21X1_509 ( .gnd(gnd), .vdd(vdd), .A(_5309_), .B(_4547__bF_buf61), .C(_5310_), .Y(_3677__2_) );
INVX1 INVX1_443 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__3_), .Y(_5311_) );
AOI22X1 AOI22X1_547 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf58), .B(block[35]), .C(w_mem_inst_w_mem_14__3_), .D(_4548__bF_buf60), .Y(_5312_) );
OAI21X1 OAI21X1_510 ( .gnd(gnd), .vdd(vdd), .A(_5311_), .B(_4547__bF_buf60), .C(_5312_), .Y(_3677__3_) );
INVX1 INVX1_444 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__4_), .Y(_5313_) );
AOI22X1 AOI22X1_548 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf57), .B(block[36]), .C(w_mem_inst_w_mem_14__4_), .D(_4548__bF_buf59), .Y(_5314_) );
OAI21X1 OAI21X1_511 ( .gnd(gnd), .vdd(vdd), .A(_5313_), .B(_4547__bF_buf59), .C(_5314_), .Y(_3677__4_) );
INVX1 INVX1_445 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__5_), .Y(_5315_) );
AOI22X1 AOI22X1_549 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf56), .B(block[37]), .C(w_mem_inst_w_mem_14__5_), .D(_4548__bF_buf58), .Y(_5316_) );
OAI21X1 OAI21X1_512 ( .gnd(gnd), .vdd(vdd), .A(_5315_), .B(_4547__bF_buf58), .C(_5316_), .Y(_3677__5_) );
INVX1 INVX1_446 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__6_), .Y(_5317_) );
AOI22X1 AOI22X1_550 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf55), .B(block[38]), .C(w_mem_inst_w_mem_14__6_), .D(_4548__bF_buf57), .Y(_5318_) );
OAI21X1 OAI21X1_513 ( .gnd(gnd), .vdd(vdd), .A(_5317_), .B(_4547__bF_buf57), .C(_5318_), .Y(_3677__6_) );
INVX1 INVX1_447 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__7_), .Y(_5319_) );
AOI22X1 AOI22X1_551 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf54), .B(block[39]), .C(w_mem_inst_w_mem_14__7_), .D(_4548__bF_buf56), .Y(_5320_) );
OAI21X1 OAI21X1_514 ( .gnd(gnd), .vdd(vdd), .A(_5319_), .B(_4547__bF_buf56), .C(_5320_), .Y(_3677__7_) );
INVX1 INVX1_448 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__8_), .Y(_5321_) );
AOI22X1 AOI22X1_552 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf53), .B(block[40]), .C(w_mem_inst_w_mem_14__8_), .D(_4548__bF_buf55), .Y(_5322_) );
OAI21X1 OAI21X1_515 ( .gnd(gnd), .vdd(vdd), .A(_5321_), .B(_4547__bF_buf55), .C(_5322_), .Y(_3677__8_) );
INVX1 INVX1_449 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__9_), .Y(_5323_) );
AOI22X1 AOI22X1_553 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf52), .B(block[41]), .C(w_mem_inst_w_mem_14__9_), .D(_4548__bF_buf54), .Y(_5324_) );
OAI21X1 OAI21X1_516 ( .gnd(gnd), .vdd(vdd), .A(_5323_), .B(_4547__bF_buf54), .C(_5324_), .Y(_3677__9_) );
INVX1 INVX1_450 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__10_), .Y(_5325_) );
AOI22X1 AOI22X1_554 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf51), .B(block[42]), .C(w_mem_inst_w_mem_14__10_), .D(_4548__bF_buf53), .Y(_5326_) );
OAI21X1 OAI21X1_517 ( .gnd(gnd), .vdd(vdd), .A(_5325_), .B(_4547__bF_buf53), .C(_5326_), .Y(_3677__10_) );
INVX1 INVX1_451 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__11_), .Y(_5327_) );
AOI22X1 AOI22X1_555 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf50), .B(block[43]), .C(w_mem_inst_w_mem_14__11_), .D(_4548__bF_buf52), .Y(_5328_) );
OAI21X1 OAI21X1_518 ( .gnd(gnd), .vdd(vdd), .A(_5327_), .B(_4547__bF_buf52), .C(_5328_), .Y(_3677__11_) );
INVX1 INVX1_452 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__12_), .Y(_5329_) );
AOI22X1 AOI22X1_556 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf49), .B(block[44]), .C(w_mem_inst_w_mem_14__12_), .D(_4548__bF_buf51), .Y(_5330_) );
OAI21X1 OAI21X1_519 ( .gnd(gnd), .vdd(vdd), .A(_5329_), .B(_4547__bF_buf51), .C(_5330_), .Y(_3677__12_) );
INVX1 INVX1_453 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__13_), .Y(_5331_) );
AOI22X1 AOI22X1_557 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf48), .B(block[45]), .C(w_mem_inst_w_mem_14__13_), .D(_4548__bF_buf50), .Y(_5332_) );
OAI21X1 OAI21X1_520 ( .gnd(gnd), .vdd(vdd), .A(_5331_), .B(_4547__bF_buf50), .C(_5332_), .Y(_3677__13_) );
INVX1 INVX1_454 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__14_), .Y(_5333_) );
AOI22X1 AOI22X1_558 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf47), .B(block[46]), .C(w_mem_inst_w_mem_14__14_), .D(_4548__bF_buf49), .Y(_5334_) );
OAI21X1 OAI21X1_521 ( .gnd(gnd), .vdd(vdd), .A(_5333_), .B(_4547__bF_buf49), .C(_5334_), .Y(_3677__14_) );
INVX1 INVX1_455 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__15_), .Y(_5335_) );
AOI22X1 AOI22X1_559 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf46), .B(block[47]), .C(w_mem_inst_w_mem_14__15_), .D(_4548__bF_buf48), .Y(_5336_) );
OAI21X1 OAI21X1_522 ( .gnd(gnd), .vdd(vdd), .A(_5335_), .B(_4547__bF_buf48), .C(_5336_), .Y(_3677__15_) );
INVX1 INVX1_456 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__16_), .Y(_5337_) );
AOI22X1 AOI22X1_560 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf45), .B(block[48]), .C(w_mem_inst_w_mem_14__16_), .D(_4548__bF_buf47), .Y(_5338_) );
OAI21X1 OAI21X1_523 ( .gnd(gnd), .vdd(vdd), .A(_5337_), .B(_4547__bF_buf47), .C(_5338_), .Y(_3677__16_) );
INVX1 INVX1_457 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__17_), .Y(_5339_) );
AOI22X1 AOI22X1_561 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf44), .B(block[49]), .C(w_mem_inst_w_mem_14__17_), .D(_4548__bF_buf46), .Y(_5340_) );
OAI21X1 OAI21X1_524 ( .gnd(gnd), .vdd(vdd), .A(_5339_), .B(_4547__bF_buf46), .C(_5340_), .Y(_3677__17_) );
INVX1 INVX1_458 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__18_), .Y(_5341_) );
AOI22X1 AOI22X1_562 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf43), .B(block[50]), .C(w_mem_inst_w_mem_14__18_), .D(_4548__bF_buf45), .Y(_5342_) );
OAI21X1 OAI21X1_525 ( .gnd(gnd), .vdd(vdd), .A(_5341_), .B(_4547__bF_buf45), .C(_5342_), .Y(_3677__18_) );
INVX1 INVX1_459 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__19_), .Y(_5343_) );
AOI22X1 AOI22X1_563 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf42), .B(block[51]), .C(w_mem_inst_w_mem_14__19_), .D(_4548__bF_buf44), .Y(_5344_) );
OAI21X1 OAI21X1_526 ( .gnd(gnd), .vdd(vdd), .A(_5343_), .B(_4547__bF_buf44), .C(_5344_), .Y(_3677__19_) );
INVX1 INVX1_460 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__20_), .Y(_5345_) );
AOI22X1 AOI22X1_564 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf41), .B(block[52]), .C(w_mem_inst_w_mem_14__20_), .D(_4548__bF_buf43), .Y(_5346_) );
OAI21X1 OAI21X1_527 ( .gnd(gnd), .vdd(vdd), .A(_5345_), .B(_4547__bF_buf43), .C(_5346_), .Y(_3677__20_) );
INVX1 INVX1_461 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__21_), .Y(_5347_) );
AOI22X1 AOI22X1_565 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf40), .B(block[53]), .C(w_mem_inst_w_mem_14__21_), .D(_4548__bF_buf42), .Y(_5348_) );
OAI21X1 OAI21X1_528 ( .gnd(gnd), .vdd(vdd), .A(_5347_), .B(_4547__bF_buf42), .C(_5348_), .Y(_3677__21_) );
INVX1 INVX1_462 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__22_), .Y(_5349_) );
AOI22X1 AOI22X1_566 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf39), .B(block[54]), .C(w_mem_inst_w_mem_14__22_), .D(_4548__bF_buf41), .Y(_5350_) );
OAI21X1 OAI21X1_529 ( .gnd(gnd), .vdd(vdd), .A(_5349_), .B(_4547__bF_buf41), .C(_5350_), .Y(_3677__22_) );
INVX1 INVX1_463 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__23_), .Y(_5351_) );
AOI22X1 AOI22X1_567 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf38), .B(block[55]), .C(w_mem_inst_w_mem_14__23_), .D(_4548__bF_buf40), .Y(_5352_) );
OAI21X1 OAI21X1_530 ( .gnd(gnd), .vdd(vdd), .A(_5351_), .B(_4547__bF_buf40), .C(_5352_), .Y(_3677__23_) );
INVX1 INVX1_464 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__24_), .Y(_5353_) );
AOI22X1 AOI22X1_568 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf37), .B(block[56]), .C(w_mem_inst_w_mem_14__24_), .D(_4548__bF_buf39), .Y(_5354_) );
OAI21X1 OAI21X1_531 ( .gnd(gnd), .vdd(vdd), .A(_5353_), .B(_4547__bF_buf39), .C(_5354_), .Y(_3677__24_) );
INVX1 INVX1_465 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__25_), .Y(_5355_) );
AOI22X1 AOI22X1_569 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf36), .B(block[57]), .C(w_mem_inst_w_mem_14__25_), .D(_4548__bF_buf38), .Y(_5356_) );
OAI21X1 OAI21X1_532 ( .gnd(gnd), .vdd(vdd), .A(_5355_), .B(_4547__bF_buf38), .C(_5356_), .Y(_3677__25_) );
INVX1 INVX1_466 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__26_), .Y(_5357_) );
AOI22X1 AOI22X1_570 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf35), .B(block[58]), .C(w_mem_inst_w_mem_14__26_), .D(_4548__bF_buf37), .Y(_5358_) );
OAI21X1 OAI21X1_533 ( .gnd(gnd), .vdd(vdd), .A(_5357_), .B(_4547__bF_buf37), .C(_5358_), .Y(_3677__26_) );
INVX1 INVX1_467 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__27_), .Y(_5359_) );
AOI22X1 AOI22X1_571 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf34), .B(block[59]), .C(w_mem_inst_w_mem_14__27_), .D(_4548__bF_buf36), .Y(_5360_) );
OAI21X1 OAI21X1_534 ( .gnd(gnd), .vdd(vdd), .A(_5359_), .B(_4547__bF_buf36), .C(_5360_), .Y(_3677__27_) );
INVX1 INVX1_468 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__28_), .Y(_5361_) );
AOI22X1 AOI22X1_572 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf33), .B(block[60]), .C(w_mem_inst_w_mem_14__28_), .D(_4548__bF_buf35), .Y(_5362_) );
OAI21X1 OAI21X1_535 ( .gnd(gnd), .vdd(vdd), .A(_5361_), .B(_4547__bF_buf35), .C(_5362_), .Y(_3677__28_) );
INVX1 INVX1_469 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__29_), .Y(_5363_) );
AOI22X1 AOI22X1_573 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf32), .B(block[61]), .C(w_mem_inst_w_mem_14__29_), .D(_4548__bF_buf34), .Y(_5364_) );
OAI21X1 OAI21X1_536 ( .gnd(gnd), .vdd(vdd), .A(_5363_), .B(_4547__bF_buf34), .C(_5364_), .Y(_3677__29_) );
INVX1 INVX1_470 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__30_), .Y(_5365_) );
AOI22X1 AOI22X1_574 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf31), .B(block[62]), .C(w_mem_inst_w_mem_14__30_), .D(_4548__bF_buf33), .Y(_5366_) );
OAI21X1 OAI21X1_537 ( .gnd(gnd), .vdd(vdd), .A(_5365_), .B(_4547__bF_buf33), .C(_5366_), .Y(_3677__30_) );
INVX1 INVX1_471 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__31_), .Y(_5367_) );
AOI22X1 AOI22X1_575 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf30), .B(block[63]), .C(w_mem_inst_w_mem_14__31_), .D(_4548__bF_buf32), .Y(_5368_) );
OAI21X1 OAI21X1_538 ( .gnd(gnd), .vdd(vdd), .A(_5367_), .B(_4547__bF_buf32), .C(_5368_), .Y(_3677__31_) );
AOI22X1 AOI22X1_576 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf29), .B(block[0]), .C(w_mem_inst_w_mem_15__0_), .D(_4548__bF_buf31), .Y(_5369_) );
OAI21X1 OAI21X1_539 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf31), .B(_3695_), .C(_5369_), .Y(_3678__0_) );
AOI22X1 AOI22X1_577 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf28), .B(block[1]), .C(w_mem_inst_w_mem_15__1_), .D(_4548__bF_buf30), .Y(_5370_) );
OAI21X1 OAI21X1_540 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf30), .B(_3754_), .C(_5370_), .Y(_3678__1_) );
AOI22X1 AOI22X1_578 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf27), .B(block[2]), .C(w_mem_inst_w_mem_15__2_), .D(_4548__bF_buf29), .Y(_5371_) );
OAI21X1 OAI21X1_541 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf29), .B(_3781_), .C(_5371_), .Y(_3678__2_) );
AOI22X1 AOI22X1_579 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf26), .B(block[3]), .C(w_mem_inst_w_mem_15__3_), .D(_4548__bF_buf28), .Y(_5372_) );
OAI21X1 OAI21X1_542 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf28), .B(_3807_), .C(_5372_), .Y(_3678__3_) );
AOI22X1 AOI22X1_580 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf25), .B(block[4]), .C(w_mem_inst_w_mem_15__4_), .D(_4548__bF_buf27), .Y(_5373_) );
OAI21X1 OAI21X1_543 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf27), .B(_3831_), .C(_5373_), .Y(_3678__4_) );
AOI22X1 AOI22X1_581 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf24), .B(block[5]), .C(w_mem_inst_w_mem_15__5_), .D(_4548__bF_buf26), .Y(_5374_) );
OAI21X1 OAI21X1_544 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf26), .B(_3859_), .C(_5374_), .Y(_3678__5_) );
AOI22X1 AOI22X1_582 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf23), .B(block[6]), .C(w_mem_inst_w_mem_15__6_), .D(_4548__bF_buf25), .Y(_5375_) );
OAI21X1 OAI21X1_545 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf25), .B(_3884_), .C(_5375_), .Y(_3678__6_) );
AOI22X1 AOI22X1_583 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf22), .B(block[7]), .C(w_mem_inst_w_mem_15__7_), .D(_4548__bF_buf24), .Y(_5376_) );
OAI21X1 OAI21X1_546 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf24), .B(_3908_), .C(_5376_), .Y(_3678__7_) );
AOI22X1 AOI22X1_584 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf21), .B(block[8]), .C(w_mem_inst_w_mem_15__8_), .D(_4548__bF_buf23), .Y(_5377_) );
OAI21X1 OAI21X1_547 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf23), .B(_3932_), .C(_5377_), .Y(_3678__8_) );
AOI22X1 AOI22X1_585 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf20), .B(block[9]), .C(w_mem_inst_w_mem_15__9_), .D(_4548__bF_buf22), .Y(_5378_) );
OAI21X1 OAI21X1_548 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf22), .B(_3957_), .C(_5378_), .Y(_3678__9_) );
AOI22X1 AOI22X1_586 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf19), .B(block[10]), .C(w_mem_inst_w_mem_15__10_), .D(_4548__bF_buf21), .Y(_5379_) );
OAI21X1 OAI21X1_549 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf21), .B(_3982_), .C(_5379_), .Y(_3678__10_) );
AOI22X1 AOI22X1_587 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf18), .B(block[11]), .C(w_mem_inst_w_mem_15__11_), .D(_4548__bF_buf20), .Y(_5380_) );
OAI21X1 OAI21X1_550 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf20), .B(_4007_), .C(_5380_), .Y(_3678__11_) );
AOI22X1 AOI22X1_588 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf17), .B(block[12]), .C(w_mem_inst_w_mem_15__12_), .D(_4548__bF_buf19), .Y(_5381_) );
OAI21X1 OAI21X1_551 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf19), .B(_4032_), .C(_5381_), .Y(_3678__12_) );
AOI22X1 AOI22X1_589 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf16), .B(block[13]), .C(w_mem_inst_w_mem_15__13_), .D(_4548__bF_buf18), .Y(_5382_) );
OAI21X1 OAI21X1_552 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf18), .B(_4057_), .C(_5382_), .Y(_3678__13_) );
AOI22X1 AOI22X1_590 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf15), .B(block[14]), .C(w_mem_inst_w_mem_15__14_), .D(_4548__bF_buf17), .Y(_5383_) );
OAI21X1 OAI21X1_553 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf17), .B(_4082_), .C(_5383_), .Y(_3678__14_) );
AOI22X1 AOI22X1_591 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf14), .B(block[15]), .C(w_mem_inst_w_mem_15__15_), .D(_4548__bF_buf16), .Y(_5384_) );
OAI21X1 OAI21X1_554 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf16), .B(_4106_), .C(_5384_), .Y(_3678__15_) );
AOI22X1 AOI22X1_592 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf13), .B(block[16]), .C(w_mem_inst_w_mem_15__16_), .D(_4548__bF_buf15), .Y(_5385_) );
OAI21X1 OAI21X1_555 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf15), .B(_4130_), .C(_5385_), .Y(_3678__16_) );
AOI22X1 AOI22X1_593 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf12), .B(block[17]), .C(w_mem_inst_w_mem_15__17_), .D(_4548__bF_buf14), .Y(_5386_) );
OAI21X1 OAI21X1_556 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf14), .B(_4155_), .C(_5386_), .Y(_3678__17_) );
AOI22X1 AOI22X1_594 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf11), .B(block[18]), .C(w_mem_inst_w_mem_15__18_), .D(_4548__bF_buf13), .Y(_5387_) );
OAI21X1 OAI21X1_557 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf13), .B(_4180_), .C(_5387_), .Y(_3678__18_) );
AOI22X1 AOI22X1_595 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf10), .B(block[19]), .C(w_mem_inst_w_mem_15__19_), .D(_4548__bF_buf12), .Y(_5388_) );
OAI21X1 OAI21X1_558 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf12), .B(_4205_), .C(_5388_), .Y(_3678__19_) );
AOI22X1 AOI22X1_596 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf9), .B(block[20]), .C(w_mem_inst_w_mem_15__20_), .D(_4548__bF_buf11), .Y(_5389_) );
OAI21X1 OAI21X1_559 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf11), .B(_4230_), .C(_5389_), .Y(_3678__20_) );
AOI22X1 AOI22X1_597 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf8), .B(block[21]), .C(w_mem_inst_w_mem_15__21_), .D(_4548__bF_buf10), .Y(_5390_) );
OAI21X1 OAI21X1_560 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf10), .B(_4255_), .C(_5390_), .Y(_3678__21_) );
AOI22X1 AOI22X1_598 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf7), .B(block[22]), .C(w_mem_inst_w_mem_15__22_), .D(_4548__bF_buf9), .Y(_5391_) );
OAI21X1 OAI21X1_561 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf9), .B(_4280_), .C(_5391_), .Y(_3678__22_) );
AOI22X1 AOI22X1_599 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf6), .B(block[23]), .C(w_mem_inst_w_mem_15__23_), .D(_4548__bF_buf8), .Y(_5392_) );
OAI21X1 OAI21X1_562 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf8), .B(_4304_), .C(_5392_), .Y(_3678__23_) );
AOI22X1 AOI22X1_600 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf5), .B(block[24]), .C(w_mem_inst_w_mem_15__24_), .D(_4548__bF_buf7), .Y(_5393_) );
OAI21X1 OAI21X1_563 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf7), .B(_4328_), .C(_5393_), .Y(_3678__24_) );
AOI22X1 AOI22X1_601 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf4), .B(block[25]), .C(w_mem_inst_w_mem_15__25_), .D(_4548__bF_buf6), .Y(_5394_) );
OAI21X1 OAI21X1_564 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf6), .B(_4353_), .C(_5394_), .Y(_3678__25_) );
AOI22X1 AOI22X1_602 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf3), .B(block[26]), .C(w_mem_inst_w_mem_15__26_), .D(_4548__bF_buf5), .Y(_5395_) );
OAI21X1 OAI21X1_565 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf5), .B(_4378_), .C(_5395_), .Y(_3678__26_) );
AOI22X1 AOI22X1_603 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf2), .B(block[27]), .C(w_mem_inst_w_mem_15__27_), .D(_4548__bF_buf4), .Y(_5396_) );
OAI21X1 OAI21X1_566 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf4), .B(_4403_), .C(_5396_), .Y(_3678__27_) );
AOI22X1 AOI22X1_604 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf1), .B(block[28]), .C(w_mem_inst_w_mem_15__28_), .D(_4548__bF_buf3), .Y(_5397_) );
OAI21X1 OAI21X1_567 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf3), .B(_4428_), .C(_5397_), .Y(_3678__28_) );
AOI22X1 AOI22X1_605 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf0), .B(block[29]), .C(w_mem_inst_w_mem_15__29_), .D(_4548__bF_buf2), .Y(_5398_) );
OAI21X1 OAI21X1_568 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf2), .B(_4453_), .C(_5398_), .Y(_3678__29_) );
AOI22X1 AOI22X1_606 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf63), .B(block[30]), .C(w_mem_inst_w_mem_15__30_), .D(_4548__bF_buf1), .Y(_5399_) );
OAI21X1 OAI21X1_569 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf1), .B(_4478_), .C(_5399_), .Y(_3678__30_) );
AOI22X1 AOI22X1_607 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_rst_bF_buf62), .B(block[31]), .C(w_mem_inst_w_mem_15__31_), .D(_4548__bF_buf0), .Y(_5400_) );
OAI21X1 OAI21X1_570 ( .gnd(gnd), .vdd(vdd), .A(_4547__bF_buf0), .B(_4502_), .C(_5400_), .Y(_3678__31_) );
DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_3671__0_), .Q(w_mem_inst_w_ctr_reg_0_) );
DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_3671__1_), .Q(w_mem_inst_w_ctr_reg_1_) );
DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_3671__2_), .Q(w_mem_inst_w_ctr_reg_2_) );
DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_3671__3_), .Q(w_mem_inst_w_ctr_reg_3_) );
DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_3671__4_), .Q(w_mem_inst_w_ctr_reg_4_) );
DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_3671__5_), .Q(w_mem_inst_w_ctr_reg_5_) );
DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_3671__6_), .Q(w_mem_inst_w_ctr_reg_6_) );
DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_3670_), .Q(w_mem_inst_sha1_w_mem_ctrl_reg), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_3672__0_), .Q(w_mem_inst_w_mem_0__0_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_3672__1_), .Q(w_mem_inst_w_mem_0__1_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_3672__2_), .Q(w_mem_inst_w_mem_0__2_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_3672__3_), .Q(w_mem_inst_w_mem_0__3_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_3672__4_), .Q(w_mem_inst_w_mem_0__4_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_3672__5_), .Q(w_mem_inst_w_mem_0__5_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_3672__6_), .Q(w_mem_inst_w_mem_0__6_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_3672__7_), .Q(w_mem_inst_w_mem_0__7_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_3672__8_), .Q(w_mem_inst_w_mem_0__8_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_3672__9_), .Q(w_mem_inst_w_mem_0__9_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_3672__10_), .Q(w_mem_inst_w_mem_0__10_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_3672__11_), .Q(w_mem_inst_w_mem_0__11_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_3672__12_), .Q(w_mem_inst_w_mem_0__12_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_3672__13_), .Q(w_mem_inst_w_mem_0__13_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_3672__14_), .Q(w_mem_inst_w_mem_0__14_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_3672__15_), .Q(w_mem_inst_w_mem_0__15_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_3672__16_), .Q(w_mem_inst_w_mem_0__16_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_3672__17_), .Q(w_mem_inst_w_mem_0__17_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_3672__18_), .Q(w_mem_inst_w_mem_0__18_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_3672__19_), .Q(w_mem_inst_w_mem_0__19_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_3672__20_), .Q(w_mem_inst_w_mem_0__20_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_3672__21_), .Q(w_mem_inst_w_mem_0__21_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_3672__22_), .Q(w_mem_inst_w_mem_0__22_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_3672__23_), .Q(w_mem_inst_w_mem_0__23_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_3672__24_), .Q(w_mem_inst_w_mem_0__24_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_3672__25_), .Q(w_mem_inst_w_mem_0__25_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_3672__26_), .Q(w_mem_inst_w_mem_0__26_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_3672__27_), .Q(w_mem_inst_w_mem_0__27_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_3672__28_), .Q(w_mem_inst_w_mem_0__28_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_3672__29_), .Q(w_mem_inst_w_mem_0__29_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_3672__30_), .Q(w_mem_inst_w_mem_0__30_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_3672__31_), .Q(w_mem_inst_w_mem_0__31_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_3679__0_), .Q(w_mem_inst_w_mem_1__0_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_3679__1_), .Q(w_mem_inst_w_mem_1__1_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_3679__2_), .Q(w_mem_inst_w_mem_1__2_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_3679__3_), .Q(w_mem_inst_w_mem_1__3_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_3679__4_), .Q(w_mem_inst_w_mem_1__4_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_3679__5_), .Q(w_mem_inst_w_mem_1__5_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_3679__6_), .Q(w_mem_inst_w_mem_1__6_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_3679__7_), .Q(w_mem_inst_w_mem_1__7_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_3679__8_), .Q(w_mem_inst_w_mem_1__8_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_3679__9_), .Q(w_mem_inst_w_mem_1__9_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_3679__10_), .Q(w_mem_inst_w_mem_1__10_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_3679__11_), .Q(w_mem_inst_w_mem_1__11_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_3679__12_), .Q(w_mem_inst_w_mem_1__12_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_3679__13_), .Q(w_mem_inst_w_mem_1__13_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_3679__14_), .Q(w_mem_inst_w_mem_1__14_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_3679__15_), .Q(w_mem_inst_w_mem_1__15_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_3679__16_), .Q(w_mem_inst_w_mem_1__16_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_3679__17_), .Q(w_mem_inst_w_mem_1__17_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_3679__18_), .Q(w_mem_inst_w_mem_1__18_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_3679__19_), .Q(w_mem_inst_w_mem_1__19_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_3679__20_), .Q(w_mem_inst_w_mem_1__20_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_3679__21_), .Q(w_mem_inst_w_mem_1__21_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_3679__22_), .Q(w_mem_inst_w_mem_1__22_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_3679__23_), .Q(w_mem_inst_w_mem_1__23_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_3679__24_), .Q(w_mem_inst_w_mem_1__24_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_3679__25_), .Q(w_mem_inst_w_mem_1__25_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_3679__26_), .Q(w_mem_inst_w_mem_1__26_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_3679__27_), .Q(w_mem_inst_w_mem_1__27_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_3679__28_), .Q(w_mem_inst_w_mem_1__28_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_3679__29_), .Q(w_mem_inst_w_mem_1__29_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_3679__30_), .Q(w_mem_inst_w_mem_1__30_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_3679__31_), .Q(w_mem_inst_w_mem_1__31_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_3680__0_), .Q(w_mem_inst_w_mem_2__0_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_3680__1_), .Q(w_mem_inst_w_mem_2__1_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_3680__2_), .Q(w_mem_inst_w_mem_2__2_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_3680__3_), .Q(w_mem_inst_w_mem_2__3_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_3680__4_), .Q(w_mem_inst_w_mem_2__4_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3680__5_), .Q(w_mem_inst_w_mem_2__5_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3680__6_), .Q(w_mem_inst_w_mem_2__6_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3680__7_), .Q(w_mem_inst_w_mem_2__7_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_3680__8_), .Q(w_mem_inst_w_mem_2__8_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3680__9_), .Q(w_mem_inst_w_mem_2__9_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_3680__10_), .Q(w_mem_inst_w_mem_2__10_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3680__11_), .Q(w_mem_inst_w_mem_2__11_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3680__12_), .Q(w_mem_inst_w_mem_2__12_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3680__13_), .Q(w_mem_inst_w_mem_2__13_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3680__14_), .Q(w_mem_inst_w_mem_2__14_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3680__15_), .Q(w_mem_inst_w_mem_2__15_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3680__16_), .Q(w_mem_inst_w_mem_2__16_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_3680__17_), .Q(w_mem_inst_w_mem_2__17_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_3680__18_), .Q(w_mem_inst_w_mem_2__18_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_3680__19_), .Q(w_mem_inst_w_mem_2__19_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_3680__20_), .Q(w_mem_inst_w_mem_2__20_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_3680__21_), .Q(w_mem_inst_w_mem_2__21_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_3680__22_), .Q(w_mem_inst_w_mem_2__22_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_3680__23_), .Q(w_mem_inst_w_mem_2__23_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_3680__24_), .Q(w_mem_inst_w_mem_2__24_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_3680__25_), .Q(w_mem_inst_w_mem_2__25_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_3680__26_), .Q(w_mem_inst_w_mem_2__26_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_3680__27_), .Q(w_mem_inst_w_mem_2__27_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_3680__28_), .Q(w_mem_inst_w_mem_2__28_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_3680__29_), .Q(w_mem_inst_w_mem_2__29_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_3680__30_), .Q(w_mem_inst_w_mem_2__30_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_3680__31_), .Q(w_mem_inst_w_mem_2__31_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_3681__0_), .Q(w_mem_inst_w_mem_3__0_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_3681__1_), .Q(w_mem_inst_w_mem_3__1_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_3681__2_), .Q(w_mem_inst_w_mem_3__2_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_3681__3_), .Q(w_mem_inst_w_mem_3__3_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_3681__4_), .Q(w_mem_inst_w_mem_3__4_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_3681__5_), .Q(w_mem_inst_w_mem_3__5_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_3681__6_), .Q(w_mem_inst_w_mem_3__6_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_3681__7_), .Q(w_mem_inst_w_mem_3__7_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_3681__8_), .Q(w_mem_inst_w_mem_3__8_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_3681__9_), .Q(w_mem_inst_w_mem_3__9_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_3681__10_), .Q(w_mem_inst_w_mem_3__10_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_3681__11_), .Q(w_mem_inst_w_mem_3__11_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_3681__12_), .Q(w_mem_inst_w_mem_3__12_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_3681__13_), .Q(w_mem_inst_w_mem_3__13_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_3681__14_), .Q(w_mem_inst_w_mem_3__14_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_3681__15_), .Q(w_mem_inst_w_mem_3__15_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_3681__16_), .Q(w_mem_inst_w_mem_3__16_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_3681__17_), .Q(w_mem_inst_w_mem_3__17_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_3681__18_), .Q(w_mem_inst_w_mem_3__18_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_3681__19_), .Q(w_mem_inst_w_mem_3__19_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_3681__20_), .Q(w_mem_inst_w_mem_3__20_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_3681__21_), .Q(w_mem_inst_w_mem_3__21_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_3681__22_), .Q(w_mem_inst_w_mem_3__22_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_3681__23_), .Q(w_mem_inst_w_mem_3__23_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_3681__24_), .Q(w_mem_inst_w_mem_3__24_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_3681__25_), .Q(w_mem_inst_w_mem_3__25_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_3681__26_), .Q(w_mem_inst_w_mem_3__26_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_3681__27_), .Q(w_mem_inst_w_mem_3__27_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_3681__28_), .Q(w_mem_inst_w_mem_3__28_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_3681__29_), .Q(w_mem_inst_w_mem_3__29_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_3681__30_), .Q(w_mem_inst_w_mem_3__30_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_3681__31_), .Q(w_mem_inst_w_mem_3__31_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_3682__0_), .Q(w_mem_inst_w_mem_4__0_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_3682__1_), .Q(w_mem_inst_w_mem_4__1_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_3682__2_), .Q(w_mem_inst_w_mem_4__2_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_3682__3_), .Q(w_mem_inst_w_mem_4__3_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_3682__4_), .Q(w_mem_inst_w_mem_4__4_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_3682__5_), .Q(w_mem_inst_w_mem_4__5_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_3682__6_), .Q(w_mem_inst_w_mem_4__6_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_3682__7_), .Q(w_mem_inst_w_mem_4__7_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_3682__8_), .Q(w_mem_inst_w_mem_4__8_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_3682__9_), .Q(w_mem_inst_w_mem_4__9_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_3682__10_), .Q(w_mem_inst_w_mem_4__10_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_3682__11_), .Q(w_mem_inst_w_mem_4__11_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_3682__12_), .Q(w_mem_inst_w_mem_4__12_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_3682__13_), .Q(w_mem_inst_w_mem_4__13_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_3682__14_), .Q(w_mem_inst_w_mem_4__14_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_3682__15_), .Q(w_mem_inst_w_mem_4__15_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_3682__16_), .Q(w_mem_inst_w_mem_4__16_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_3682__17_), .Q(w_mem_inst_w_mem_4__17_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_3682__18_), .Q(w_mem_inst_w_mem_4__18_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_3682__19_), .Q(w_mem_inst_w_mem_4__19_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_3682__20_), .Q(w_mem_inst_w_mem_4__20_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_3682__21_), .Q(w_mem_inst_w_mem_4__21_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_3682__22_), .Q(w_mem_inst_w_mem_4__22_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_3682__23_), .Q(w_mem_inst_w_mem_4__23_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_3682__24_), .Q(w_mem_inst_w_mem_4__24_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_3682__25_), .Q(w_mem_inst_w_mem_4__25_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_3682__26_), .Q(w_mem_inst_w_mem_4__26_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_3682__27_), .Q(w_mem_inst_w_mem_4__27_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_3682__28_), .Q(w_mem_inst_w_mem_4__28_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_3682__29_), .Q(w_mem_inst_w_mem_4__29_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3682__30_), .Q(w_mem_inst_w_mem_4__30_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3682__31_), .Q(w_mem_inst_w_mem_4__31_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3683__0_), .Q(w_mem_inst_w_mem_5__0_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_3683__1_), .Q(w_mem_inst_w_mem_5__1_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3683__2_), .Q(w_mem_inst_w_mem_5__2_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_3683__3_), .Q(w_mem_inst_w_mem_5__3_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3683__4_), .Q(w_mem_inst_w_mem_5__4_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3683__5_), .Q(w_mem_inst_w_mem_5__5_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3683__6_), .Q(w_mem_inst_w_mem_5__6_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3683__7_), .Q(w_mem_inst_w_mem_5__7_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3683__8_), .Q(w_mem_inst_w_mem_5__8_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3683__9_), .Q(w_mem_inst_w_mem_5__9_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_3683__10_), .Q(w_mem_inst_w_mem_5__10_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_3683__11_), .Q(w_mem_inst_w_mem_5__11_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_3683__12_), .Q(w_mem_inst_w_mem_5__12_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_3683__13_), .Q(w_mem_inst_w_mem_5__13_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_3683__14_), .Q(w_mem_inst_w_mem_5__14_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_3683__15_), .Q(w_mem_inst_w_mem_5__15_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_3683__16_), .Q(w_mem_inst_w_mem_5__16_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_3683__17_), .Q(w_mem_inst_w_mem_5__17_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_3683__18_), .Q(w_mem_inst_w_mem_5__18_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_3683__19_), .Q(w_mem_inst_w_mem_5__19_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_3683__20_), .Q(w_mem_inst_w_mem_5__20_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_3683__21_), .Q(w_mem_inst_w_mem_5__21_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_3683__22_), .Q(w_mem_inst_w_mem_5__22_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_3683__23_), .Q(w_mem_inst_w_mem_5__23_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_3683__24_), .Q(w_mem_inst_w_mem_5__24_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_3683__25_), .Q(w_mem_inst_w_mem_5__25_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_3683__26_), .Q(w_mem_inst_w_mem_5__26_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_3683__27_), .Q(w_mem_inst_w_mem_5__27_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_3683__28_), .Q(w_mem_inst_w_mem_5__28_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_3683__29_), .Q(w_mem_inst_w_mem_5__29_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_3683__30_), .Q(w_mem_inst_w_mem_5__30_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_3683__31_), .Q(w_mem_inst_w_mem_5__31_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_3684__0_), .Q(w_mem_inst_w_mem_6__0_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_3684__1_), .Q(w_mem_inst_w_mem_6__1_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_3684__2_), .Q(w_mem_inst_w_mem_6__2_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_3684__3_), .Q(w_mem_inst_w_mem_6__3_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_3684__4_), .Q(w_mem_inst_w_mem_6__4_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_3684__5_), .Q(w_mem_inst_w_mem_6__5_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_3684__6_), .Q(w_mem_inst_w_mem_6__6_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_3684__7_), .Q(w_mem_inst_w_mem_6__7_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_3684__8_), .Q(w_mem_inst_w_mem_6__8_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_3684__9_), .Q(w_mem_inst_w_mem_6__9_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_3684__10_), .Q(w_mem_inst_w_mem_6__10_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_3684__11_), .Q(w_mem_inst_w_mem_6__11_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_3684__12_), .Q(w_mem_inst_w_mem_6__12_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_3684__13_), .Q(w_mem_inst_w_mem_6__13_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_3684__14_), .Q(w_mem_inst_w_mem_6__14_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_3684__15_), .Q(w_mem_inst_w_mem_6__15_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_3684__16_), .Q(w_mem_inst_w_mem_6__16_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_3684__17_), .Q(w_mem_inst_w_mem_6__17_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_3684__18_), .Q(w_mem_inst_w_mem_6__18_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_3684__19_), .Q(w_mem_inst_w_mem_6__19_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_3684__20_), .Q(w_mem_inst_w_mem_6__20_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_3684__21_), .Q(w_mem_inst_w_mem_6__21_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_3684__22_), .Q(w_mem_inst_w_mem_6__22_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_3684__23_), .Q(w_mem_inst_w_mem_6__23_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_3684__24_), .Q(w_mem_inst_w_mem_6__24_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_3684__25_), .Q(w_mem_inst_w_mem_6__25_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_3684__26_), .Q(w_mem_inst_w_mem_6__26_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_3684__27_), .Q(w_mem_inst_w_mem_6__27_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_3684__28_), .Q(w_mem_inst_w_mem_6__28_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_3684__29_), .Q(w_mem_inst_w_mem_6__29_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_3684__30_), .Q(w_mem_inst_w_mem_6__30_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_3684__31_), .Q(w_mem_inst_w_mem_6__31_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_3685__0_), .Q(w_mem_inst_w_mem_7__0_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_3685__1_), .Q(w_mem_inst_w_mem_7__1_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_3685__2_), .Q(w_mem_inst_w_mem_7__2_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_3685__3_), .Q(w_mem_inst_w_mem_7__3_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_3685__4_), .Q(w_mem_inst_w_mem_7__4_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_3685__5_), .Q(w_mem_inst_w_mem_7__5_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_3685__6_), .Q(w_mem_inst_w_mem_7__6_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_3685__7_), .Q(w_mem_inst_w_mem_7__7_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_3685__8_), .Q(w_mem_inst_w_mem_7__8_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_3685__9_), .Q(w_mem_inst_w_mem_7__9_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_3685__10_), .Q(w_mem_inst_w_mem_7__10_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_3685__11_), .Q(w_mem_inst_w_mem_7__11_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_3685__12_), .Q(w_mem_inst_w_mem_7__12_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_3685__13_), .Q(w_mem_inst_w_mem_7__13_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_3685__14_), .Q(w_mem_inst_w_mem_7__14_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_3685__15_), .Q(w_mem_inst_w_mem_7__15_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_3685__16_), .Q(w_mem_inst_w_mem_7__16_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_3685__17_), .Q(w_mem_inst_w_mem_7__17_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_3685__18_), .Q(w_mem_inst_w_mem_7__18_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_3685__19_), .Q(w_mem_inst_w_mem_7__19_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_3685__20_), .Q(w_mem_inst_w_mem_7__20_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_3685__21_), .Q(w_mem_inst_w_mem_7__21_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_3685__22_), .Q(w_mem_inst_w_mem_7__22_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3685__23_), .Q(w_mem_inst_w_mem_7__23_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3685__24_), .Q(w_mem_inst_w_mem_7__24_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3685__25_), .Q(w_mem_inst_w_mem_7__25_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_3685__26_), .Q(w_mem_inst_w_mem_7__26_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3685__27_), .Q(w_mem_inst_w_mem_7__27_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_3685__28_), .Q(w_mem_inst_w_mem_7__28_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3685__29_), .Q(w_mem_inst_w_mem_7__29_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3685__30_), .Q(w_mem_inst_w_mem_7__30_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3685__31_), .Q(w_mem_inst_w_mem_7__31_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3686__0_), .Q(w_mem_inst_w_mem_8__0_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3686__1_), .Q(w_mem_inst_w_mem_8__1_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3686__2_), .Q(w_mem_inst_w_mem_8__2_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_3686__3_), .Q(w_mem_inst_w_mem_8__3_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_3686__4_), .Q(w_mem_inst_w_mem_8__4_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_3686__5_), .Q(w_mem_inst_w_mem_8__5_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_3686__6_), .Q(w_mem_inst_w_mem_8__6_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_3686__7_), .Q(w_mem_inst_w_mem_8__7_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_3686__8_), .Q(w_mem_inst_w_mem_8__8_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_3686__9_), .Q(w_mem_inst_w_mem_8__9_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_3686__10_), .Q(w_mem_inst_w_mem_8__10_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_3686__11_), .Q(w_mem_inst_w_mem_8__11_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_3686__12_), .Q(w_mem_inst_w_mem_8__12_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_3686__13_), .Q(w_mem_inst_w_mem_8__13_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_3686__14_), .Q(w_mem_inst_w_mem_8__14_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_3686__15_), .Q(w_mem_inst_w_mem_8__15_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_3686__16_), .Q(w_mem_inst_w_mem_8__16_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_3686__17_), .Q(w_mem_inst_w_mem_8__17_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_3686__18_), .Q(w_mem_inst_w_mem_8__18_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_3686__19_), .Q(w_mem_inst_w_mem_8__19_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_3686__20_), .Q(w_mem_inst_w_mem_8__20_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_3686__21_), .Q(w_mem_inst_w_mem_8__21_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_3686__22_), .Q(w_mem_inst_w_mem_8__22_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_3686__23_), .Q(w_mem_inst_w_mem_8__23_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_3686__24_), .Q(w_mem_inst_w_mem_8__24_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_3686__25_), .Q(w_mem_inst_w_mem_8__25_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_3686__26_), .Q(w_mem_inst_w_mem_8__26_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_3686__27_), .Q(w_mem_inst_w_mem_8__27_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_3686__28_), .Q(w_mem_inst_w_mem_8__28_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_3686__29_), .Q(w_mem_inst_w_mem_8__29_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_3686__30_), .Q(w_mem_inst_w_mem_8__30_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_3686__31_), .Q(w_mem_inst_w_mem_8__31_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_3687__0_), .Q(w_mem_inst_w_mem_9__0_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_3687__1_), .Q(w_mem_inst_w_mem_9__1_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_3687__2_), .Q(w_mem_inst_w_mem_9__2_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_3687__3_), .Q(w_mem_inst_w_mem_9__3_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_3687__4_), .Q(w_mem_inst_w_mem_9__4_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_3687__5_), .Q(w_mem_inst_w_mem_9__5_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_3687__6_), .Q(w_mem_inst_w_mem_9__6_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_3687__7_), .Q(w_mem_inst_w_mem_9__7_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_3687__8_), .Q(w_mem_inst_w_mem_9__8_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_3687__9_), .Q(w_mem_inst_w_mem_9__9_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_3687__10_), .Q(w_mem_inst_w_mem_9__10_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_3687__11_), .Q(w_mem_inst_w_mem_9__11_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_3687__12_), .Q(w_mem_inst_w_mem_9__12_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_3687__13_), .Q(w_mem_inst_w_mem_9__13_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_3687__14_), .Q(w_mem_inst_w_mem_9__14_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_3687__15_), .Q(w_mem_inst_w_mem_9__15_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_3687__16_), .Q(w_mem_inst_w_mem_9__16_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_3687__17_), .Q(w_mem_inst_w_mem_9__17_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_3687__18_), .Q(w_mem_inst_w_mem_9__18_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_3687__19_), .Q(w_mem_inst_w_mem_9__19_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_3687__20_), .Q(w_mem_inst_w_mem_9__20_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_3687__21_), .Q(w_mem_inst_w_mem_9__21_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_3687__22_), .Q(w_mem_inst_w_mem_9__22_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_3687__23_), .Q(w_mem_inst_w_mem_9__23_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_3687__24_), .Q(w_mem_inst_w_mem_9__24_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_3687__25_), .Q(w_mem_inst_w_mem_9__25_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_3687__26_), .Q(w_mem_inst_w_mem_9__26_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_3687__27_), .Q(w_mem_inst_w_mem_9__27_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_3687__28_), .Q(w_mem_inst_w_mem_9__28_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_3687__29_), .Q(w_mem_inst_w_mem_9__29_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_3687__30_), .Q(w_mem_inst_w_mem_9__30_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_3687__31_), .Q(w_mem_inst_w_mem_9__31_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_3673__0_), .Q(w_mem_inst_w_mem_10__0_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_3673__1_), .Q(w_mem_inst_w_mem_10__1_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_3673__2_), .Q(w_mem_inst_w_mem_10__2_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_3673__3_), .Q(w_mem_inst_w_mem_10__3_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_3673__4_), .Q(w_mem_inst_w_mem_10__4_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_3673__5_), .Q(w_mem_inst_w_mem_10__5_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_3673__6_), .Q(w_mem_inst_w_mem_10__6_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_3673__7_), .Q(w_mem_inst_w_mem_10__7_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_3673__8_), .Q(w_mem_inst_w_mem_10__8_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_3673__9_), .Q(w_mem_inst_w_mem_10__9_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_3673__10_), .Q(w_mem_inst_w_mem_10__10_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_3673__11_), .Q(w_mem_inst_w_mem_10__11_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_3673__12_), .Q(w_mem_inst_w_mem_10__12_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_3673__13_), .Q(w_mem_inst_w_mem_10__13_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_3673__14_), .Q(w_mem_inst_w_mem_10__14_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_3673__15_), .Q(w_mem_inst_w_mem_10__15_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3673__16_), .Q(w_mem_inst_w_mem_10__16_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3673__17_), .Q(w_mem_inst_w_mem_10__17_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3673__18_), .Q(w_mem_inst_w_mem_10__18_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_3673__19_), .Q(w_mem_inst_w_mem_10__19_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3673__20_), .Q(w_mem_inst_w_mem_10__20_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_3673__21_), .Q(w_mem_inst_w_mem_10__21_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3673__22_), .Q(w_mem_inst_w_mem_10__22_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3673__23_), .Q(w_mem_inst_w_mem_10__23_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3673__24_), .Q(w_mem_inst_w_mem_10__24_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3673__25_), .Q(w_mem_inst_w_mem_10__25_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3673__26_), .Q(w_mem_inst_w_mem_10__26_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3673__27_), .Q(w_mem_inst_w_mem_10__27_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_3673__28_), .Q(w_mem_inst_w_mem_10__28_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_3673__29_), .Q(w_mem_inst_w_mem_10__29_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_3673__30_), .Q(w_mem_inst_w_mem_10__30_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_3673__31_), .Q(w_mem_inst_w_mem_10__31_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_3674__0_), .Q(w_mem_inst_w_mem_11__0_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_3674__1_), .Q(w_mem_inst_w_mem_11__1_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_3674__2_), .Q(w_mem_inst_w_mem_11__2_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_3674__3_), .Q(w_mem_inst_w_mem_11__3_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_3674__4_), .Q(w_mem_inst_w_mem_11__4_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_3674__5_), .Q(w_mem_inst_w_mem_11__5_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_3674__6_), .Q(w_mem_inst_w_mem_11__6_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_3674__7_), .Q(w_mem_inst_w_mem_11__7_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_3674__8_), .Q(w_mem_inst_w_mem_11__8_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_3674__9_), .Q(w_mem_inst_w_mem_11__9_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_3674__10_), .Q(w_mem_inst_w_mem_11__10_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_3674__11_), .Q(w_mem_inst_w_mem_11__11_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_3674__12_), .Q(w_mem_inst_w_mem_11__12_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_3674__13_), .Q(w_mem_inst_w_mem_11__13_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_3674__14_), .Q(w_mem_inst_w_mem_11__14_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_3674__15_), .Q(w_mem_inst_w_mem_11__15_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_3674__16_), .Q(w_mem_inst_w_mem_11__16_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_3674__17_), .Q(w_mem_inst_w_mem_11__17_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_3674__18_), .Q(w_mem_inst_w_mem_11__18_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_3674__19_), .Q(w_mem_inst_w_mem_11__19_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_3674__20_), .Q(w_mem_inst_w_mem_11__20_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_3674__21_), .Q(w_mem_inst_w_mem_11__21_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_3674__22_), .Q(w_mem_inst_w_mem_11__22_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_3674__23_), .Q(w_mem_inst_w_mem_11__23_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_3674__24_), .Q(w_mem_inst_w_mem_11__24_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_3674__25_), .Q(w_mem_inst_w_mem_11__25_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_3674__26_), .Q(w_mem_inst_w_mem_11__26_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_3674__27_), .Q(w_mem_inst_w_mem_11__27_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_3674__28_), .Q(w_mem_inst_w_mem_11__28_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_3674__29_), .Q(w_mem_inst_w_mem_11__29_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_3674__30_), .Q(w_mem_inst_w_mem_11__30_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_3674__31_), .Q(w_mem_inst_w_mem_11__31_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_3675__0_), .Q(w_mem_inst_w_mem_12__0_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_3675__1_), .Q(w_mem_inst_w_mem_12__1_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_3675__2_), .Q(w_mem_inst_w_mem_12__2_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_3675__3_), .Q(w_mem_inst_w_mem_12__3_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_3675__4_), .Q(w_mem_inst_w_mem_12__4_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_3675__5_), .Q(w_mem_inst_w_mem_12__5_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_3675__6_), .Q(w_mem_inst_w_mem_12__6_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_3675__7_), .Q(w_mem_inst_w_mem_12__7_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_3675__8_), .Q(w_mem_inst_w_mem_12__8_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_3675__9_), .Q(w_mem_inst_w_mem_12__9_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_3675__10_), .Q(w_mem_inst_w_mem_12__10_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_3675__11_), .Q(w_mem_inst_w_mem_12__11_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_3675__12_), .Q(w_mem_inst_w_mem_12__12_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_3675__13_), .Q(w_mem_inst_w_mem_12__13_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_3675__14_), .Q(w_mem_inst_w_mem_12__14_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_3675__15_), .Q(w_mem_inst_w_mem_12__15_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_3675__16_), .Q(w_mem_inst_w_mem_12__16_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_3675__17_), .Q(w_mem_inst_w_mem_12__17_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_3675__18_), .Q(w_mem_inst_w_mem_12__18_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_3675__19_), .Q(w_mem_inst_w_mem_12__19_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_3675__20_), .Q(w_mem_inst_w_mem_12__20_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_3675__21_), .Q(w_mem_inst_w_mem_12__21_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_3675__22_), .Q(w_mem_inst_w_mem_12__22_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_3675__23_), .Q(w_mem_inst_w_mem_12__23_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_3675__24_), .Q(w_mem_inst_w_mem_12__24_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_3675__25_), .Q(w_mem_inst_w_mem_12__25_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_3675__26_), .Q(w_mem_inst_w_mem_12__26_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_3675__27_), .Q(w_mem_inst_w_mem_12__27_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_3675__28_), .Q(w_mem_inst_w_mem_12__28_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_3675__29_), .Q(w_mem_inst_w_mem_12__29_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_3675__30_), .Q(w_mem_inst_w_mem_12__30_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_3675__31_), .Q(w_mem_inst_w_mem_12__31_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_3676__0_), .Q(w_mem_inst_w_mem_13__0_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_3676__1_), .Q(w_mem_inst_w_mem_13__1_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_3676__2_), .Q(w_mem_inst_w_mem_13__2_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_3676__3_), .Q(w_mem_inst_w_mem_13__3_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_3676__4_), .Q(w_mem_inst_w_mem_13__4_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_3676__5_), .Q(w_mem_inst_w_mem_13__5_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_3676__6_), .Q(w_mem_inst_w_mem_13__6_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_3676__7_), .Q(w_mem_inst_w_mem_13__7_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_3676__8_), .Q(w_mem_inst_w_mem_13__8_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3676__9_), .Q(w_mem_inst_w_mem_13__9_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3676__10_), .Q(w_mem_inst_w_mem_13__10_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3676__11_), .Q(w_mem_inst_w_mem_13__11_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_3676__12_), .Q(w_mem_inst_w_mem_13__12_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3676__13_), .Q(w_mem_inst_w_mem_13__13_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_3676__14_), .Q(w_mem_inst_w_mem_13__14_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3676__15_), .Q(w_mem_inst_w_mem_13__15_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3676__16_), .Q(w_mem_inst_w_mem_13__16_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3676__17_), .Q(w_mem_inst_w_mem_13__17_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3676__18_), .Q(w_mem_inst_w_mem_13__18_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3676__19_), .Q(w_mem_inst_w_mem_13__19_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3676__20_), .Q(w_mem_inst_w_mem_13__20_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_3676__21_), .Q(w_mem_inst_w_mem_13__21_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_3676__22_), .Q(w_mem_inst_w_mem_13__22_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_441 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_3676__23_), .Q(w_mem_inst_w_mem_13__23_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_442 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_3676__24_), .Q(w_mem_inst_w_mem_13__24_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_443 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_3676__25_), .Q(w_mem_inst_w_mem_13__25_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_444 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_3676__26_), .Q(w_mem_inst_w_mem_13__26_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_445 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_3676__27_), .Q(w_mem_inst_w_mem_13__27_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_446 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_3676__28_), .Q(w_mem_inst_w_mem_13__28_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_447 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_3676__29_), .Q(w_mem_inst_w_mem_13__29_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_448 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_3676__30_), .Q(w_mem_inst_w_mem_13__30_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_449 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_3676__31_), .Q(w_mem_inst_w_mem_13__31_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_450 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_3677__0_), .Q(w_mem_inst_w_mem_14__0_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_451 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_3677__1_), .Q(w_mem_inst_w_mem_14__1_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_452 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_3677__2_), .Q(w_mem_inst_w_mem_14__2_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_453 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_3677__3_), .Q(w_mem_inst_w_mem_14__3_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_454 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_3677__4_), .Q(w_mem_inst_w_mem_14__4_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_455 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_3677__5_), .Q(w_mem_inst_w_mem_14__5_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_456 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_3677__6_), .Q(w_mem_inst_w_mem_14__6_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_457 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_3677__7_), .Q(w_mem_inst_w_mem_14__7_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_458 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_3677__8_), .Q(w_mem_inst_w_mem_14__8_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_459 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_3677__9_), .Q(w_mem_inst_w_mem_14__9_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_460 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_3677__10_), .Q(w_mem_inst_w_mem_14__10_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_461 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_3677__11_), .Q(w_mem_inst_w_mem_14__11_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_462 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_3677__12_), .Q(w_mem_inst_w_mem_14__12_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_463 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_3677__13_), .Q(w_mem_inst_w_mem_14__13_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_464 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_3677__14_), .Q(w_mem_inst_w_mem_14__14_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_465 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_3677__15_), .Q(w_mem_inst_w_mem_14__15_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_466 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_3677__16_), .Q(w_mem_inst_w_mem_14__16_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_467 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_3677__17_), .Q(w_mem_inst_w_mem_14__17_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_468 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_3677__18_), .Q(w_mem_inst_w_mem_14__18_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_469 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_3677__19_), .Q(w_mem_inst_w_mem_14__19_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_470 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_3677__20_), .Q(w_mem_inst_w_mem_14__20_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_471 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_3677__21_), .Q(w_mem_inst_w_mem_14__21_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_472 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_3677__22_), .Q(w_mem_inst_w_mem_14__22_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_473 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_3677__23_), .Q(w_mem_inst_w_mem_14__23_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_474 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_3677__24_), .Q(w_mem_inst_w_mem_14__24_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_475 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_3677__25_), .Q(w_mem_inst_w_mem_14__25_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_476 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_3677__26_), .Q(w_mem_inst_w_mem_14__26_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_477 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_3677__27_), .Q(w_mem_inst_w_mem_14__27_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_478 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_3677__28_), .Q(w_mem_inst_w_mem_14__28_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_479 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_3677__29_), .Q(w_mem_inst_w_mem_14__29_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_480 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_3677__30_), .Q(w_mem_inst_w_mem_14__30_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_481 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_3677__31_), .Q(w_mem_inst_w_mem_14__31_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_482 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_3678__0_), .Q(w_mem_inst_w_mem_15__0_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_483 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_3678__1_), .Q(w_mem_inst_w_mem_15__1_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_484 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_3678__2_), .Q(w_mem_inst_w_mem_15__2_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_485 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_3678__3_), .Q(w_mem_inst_w_mem_15__3_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_486 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_3678__4_), .Q(w_mem_inst_w_mem_15__4_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_487 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_3678__5_), .Q(w_mem_inst_w_mem_15__5_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_488 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_3678__6_), .Q(w_mem_inst_w_mem_15__6_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_489 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_3678__7_), .Q(w_mem_inst_w_mem_15__7_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_490 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_3678__8_), .Q(w_mem_inst_w_mem_15__8_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_491 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_3678__9_), .Q(w_mem_inst_w_mem_15__9_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_492 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_3678__10_), .Q(w_mem_inst_w_mem_15__10_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_493 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_3678__11_), .Q(w_mem_inst_w_mem_15__11_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_494 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_3678__12_), .Q(w_mem_inst_w_mem_15__12_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_495 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_3678__13_), .Q(w_mem_inst_w_mem_15__13_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_496 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_3678__14_), .Q(w_mem_inst_w_mem_15__14_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_497 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_3678__15_), .Q(w_mem_inst_w_mem_15__15_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_498 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_3678__16_), .Q(w_mem_inst_w_mem_15__16_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_499 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_3678__17_), .Q(w_mem_inst_w_mem_15__17_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_500 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_3678__18_), .Q(w_mem_inst_w_mem_15__18_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_501 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_3678__19_), .Q(w_mem_inst_w_mem_15__19_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_502 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_3678__20_), .Q(w_mem_inst_w_mem_15__20_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_503 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_3678__21_), .Q(w_mem_inst_w_mem_15__21_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_504 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_3678__22_), .Q(w_mem_inst_w_mem_15__22_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_505 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_3678__23_), .Q(w_mem_inst_w_mem_15__23_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_506 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_3678__24_), .Q(w_mem_inst_w_mem_15__24_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_507 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_3678__25_), .Q(w_mem_inst_w_mem_15__25_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_508 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_3678__26_), .Q(w_mem_inst_w_mem_15__26_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_509 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_3678__27_), .Q(w_mem_inst_w_mem_15__27_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_510 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_3678__28_), .Q(w_mem_inst_w_mem_15__28_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_511 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_3678__29_), .Q(w_mem_inst_w_mem_15__29_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_512 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_3678__30_), .Q(w_mem_inst_w_mem_15__30_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_513 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_3678__31_), .Q(w_mem_inst_w_mem_15__31_), .R(reset_n_bF_buf21), .S(vdd) );
OAI21X1 OAI21X1_571 ( .gnd(gnd), .vdd(vdd), .A(next), .B(init), .C(_3669_), .Y(_3370_) );
INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(_3370_), .Y(round_ctr_rst) );
NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(round_ctr_rst_bF_buf61), .Y(_3371_) );
NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .Y(_3372_) );
NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_6_), .B(_3372_), .Y(_3373_) );
INVX1 INVX1_472 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_1_), .Y(_3374_) );
INVX2 INVX2_3 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_0_), .Y(_3375_) );
NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_3375_), .Y(_3376_) );
INVX1 INVX1_473 ( .gnd(gnd), .vdd(vdd), .A(_3376_), .Y(_3377_) );
NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_3_), .B(round_ctr_reg_2_), .Y(_3378_) );
NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3378_), .B(_3377_), .Y(_3379_) );
INVX2 INVX2_4 ( .gnd(gnd), .vdd(vdd), .A(_3379_), .Y(_3380_) );
OAI21X1 OAI21X1_572 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_3380_), .C(round_ctr_inc_bF_buf10), .Y(_3381_) );
NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(next), .B(init), .Y(_3382_) );
AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_3382_), .B(_3669_), .C(digest_valid_new_bF_buf7), .Y(_3383_) );
OAI21X1 OAI21X1_573 ( .gnd(gnd), .vdd(vdd), .A(_3371_), .B(_3381_), .C(_3383_), .Y(_3666__0_) );
OAI21X1 OAI21X1_574 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf6), .B(_3381_), .C(_3370_), .Y(_3666__2_) );
INVX1 INVX1_474 ( .gnd(gnd), .vdd(vdd), .A(a_reg_0_), .Y(_3384_) );
INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .Y(_3385_) );
INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(_3669_), .Y(_3386_) );
OAI21X1 OAI21X1_575 ( .gnd(gnd), .vdd(vdd), .A(_3386__bF_buf7), .B(_3382_), .C(_3385_), .Y(_3387_) );
INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_6_), .Y(_3388_) );
NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .Y(_3389_) );
NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_3_), .B(round_ctr_reg_5_), .Y(_3390_) );
NAND3X1 NAND3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3389_), .C(_3390_), .Y(_3391_) );
INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .Y(_3392_) );
INVX1 INVX1_475 ( .gnd(gnd), .vdd(vdd), .A(d_reg_0_), .Y(_3393_) );
NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(c_reg_0_), .B(b_reg_0_), .Y(_3394_) );
INVX1 INVX1_476 ( .gnd(gnd), .vdd(vdd), .A(_3394_), .Y(_3395_) );
NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(c_reg_0_), .B(b_reg_0_), .Y(_3396_) );
NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3396_), .B(_3395_), .Y(_3397_) );
NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_3397_), .Y(_3398_) );
OAI21X1 OAI21X1_576 ( .gnd(gnd), .vdd(vdd), .A(_3396_), .B(_3395_), .C(d_reg_0_), .Y(_3399_) );
INVX1 INVX1_477 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_5_), .Y(_3400_) );
OAI21X1 OAI21X1_577 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_3_), .B(round_ctr_reg_2_), .C(round_ctr_reg_4_), .Y(_3401_) );
NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_3401_), .Y(_3402_) );
AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_3_), .B(round_ctr_reg_5_), .C(round_ctr_reg_6_), .Y(_3403_) );
AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_2_), .B(round_ctr_reg_4_), .C(round_ctr_reg_6_), .Y(_3404_) );
OAI21X1 OAI21X1_578 ( .gnd(gnd), .vdd(vdd), .A(_3403_), .B(_3404_), .C(_3391_), .Y(_3405_) );
OAI21X1 OAI21X1_579 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_6_), .B(_3402_), .C(_3405__bF_buf5), .Y(_3406_) );
AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_3398_), .B(_3399_), .C(_3406__bF_buf4), .Y(_3407_) );
NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_5_), .B(round_ctr_reg_6_), .Y(_3408_) );
NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_2_), .B(round_ctr_reg_4_), .Y(_3409_) );
NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_3_), .B(round_ctr_reg_4_), .Y(_3410_) );
NAND3X1 NAND3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_3409_), .B(_3410_), .C(_3408_), .Y(_3411_) );
INVX2 INVX2_5 ( .gnd(gnd), .vdd(vdd), .A(b_reg_0_), .Y(_3412_) );
INVX1 INVX1_478 ( .gnd(gnd), .vdd(vdd), .A(c_reg_0_), .Y(_3413_) );
OAI21X1 OAI21X1_580 ( .gnd(gnd), .vdd(vdd), .A(_3413_), .B(_3412_), .C(_3393_), .Y(_3414_) );
OAI21X1 OAI21X1_581 ( .gnd(gnd), .vdd(vdd), .A(c_reg_0_), .B(_3412_), .C(_3414_), .Y(_3415_) );
OAI21X1 OAI21X1_582 ( .gnd(gnd), .vdd(vdd), .A(c_reg_0_), .B(b_reg_0_), .C(_3414_), .Y(_3416_) );
OAI22X1 OAI22X1_42 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf4), .B(_3415_), .C(_3416_), .D(_3405__bF_buf4), .Y(_3417_) );
INVX1 INVX1_479 ( .gnd(gnd), .vdd(vdd), .A(w_0_), .Y(_3418_) );
NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(e_reg_0_), .B(a_reg_27_), .Y(_3419_) );
INVX1 INVX1_480 ( .gnd(gnd), .vdd(vdd), .A(_3419_), .Y(_3420_) );
NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(e_reg_0_), .B(a_reg_27_), .Y(_3421_) );
NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3421_), .B(_3420_), .Y(_3422_) );
XNOR2X1 XNOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3422_), .B(_3418_), .Y(_3423_) );
OAI21X1 OAI21X1_583 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_3407_), .C(_3423_), .Y(_3424_) );
INVX1 INVX1_481 ( .gnd(gnd), .vdd(vdd), .A(_3424_), .Y(_3425_) );
NOR3X1 NOR3X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3417_), .B(_3423_), .C(_3407_), .Y(_3426_) );
NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_3426_), .B(_3425_), .Y(_3427_) );
AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_3427_), .B(_3392_), .Y(_3428_) );
NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_3428_), .Y(_3429_) );
OAI21X1 OAI21X1_584 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3427_), .C(_3429_), .Y(_3430_) );
INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(init), .Y(_3431_) );
NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .Y(_3432_) );
NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(_3370_), .Y(_3433_) );
OAI21X1 OAI21X1_585 ( .gnd(gnd), .vdd(vdd), .A(_3667__128_), .B(_3432__bF_buf11), .C(_3433__bF_buf11), .Y(_3434_) );
AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_3430_), .B(_3434_), .Y(_3435_) );
OAI21X1 OAI21X1_586 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(_3387__bF_buf10), .C(_3435_), .Y(_5__0_) );
INVX1 INVX1_482 ( .gnd(gnd), .vdd(vdd), .A(a_reg_1_), .Y(_3436_) );
OAI21X1 OAI21X1_587 ( .gnd(gnd), .vdd(vdd), .A(_3378_), .B(_3389_), .C(_3388_), .Y(_3437_) );
NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(c_reg_1_), .B(b_reg_1_), .Y(_3438_) );
INVX2 INVX2_6 ( .gnd(gnd), .vdd(vdd), .A(c_reg_1_), .Y(_3439_) );
INVX2 INVX2_7 ( .gnd(gnd), .vdd(vdd), .A(b_reg_1_), .Y(_3440_) );
NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_3440_), .Y(_3441_) );
NAND3X1 NAND3X1_84 ( .gnd(gnd), .vdd(vdd), .A(d_reg_1_), .B(_3438_), .C(_3441_), .Y(_3442_) );
INVX2 INVX2_8 ( .gnd(gnd), .vdd(vdd), .A(d_reg_1_), .Y(_3443_) );
NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_3438_), .B(_3441_), .Y(_3444_) );
NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_3444_), .Y(_3445_) );
NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_3442_), .B(_3445_), .Y(_3446_) );
INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf3), .Y(_3447_) );
NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3390_), .Y(_3448_) );
OAI21X1 OAI21X1_588 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_3_), .B(round_ctr_reg_4_), .C(round_ctr_reg_5_), .Y(_3449_) );
NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3409_), .Y(_3450_) );
AOI22X1 AOI22X1_608 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3449_), .C(_3448_), .D(_3450_), .Y(_3451_) );
OAI21X1 OAI21X1_589 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_3440_), .C(_3443_), .Y(_3452_) );
AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_3452_), .B(_3441_), .Y(_3453_) );
OAI21X1 OAI21X1_590 ( .gnd(gnd), .vdd(vdd), .A(b_reg_1_), .B(_3443_), .C(_3438_), .Y(_3454_) );
AOI22X1 AOI22X1_609 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf4), .B(_3454_), .C(_3451__bF_buf4), .D(_3453_), .Y(_3455_) );
OAI21X1 OAI21X1_591 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf3), .B(_3446_), .C(_3455_), .Y(_3456_) );
OAI21X1 OAI21X1_592 ( .gnd(gnd), .vdd(vdd), .A(_3418_), .B(_3421_), .C(_3419_), .Y(_3457_) );
INVX1 INVX1_483 ( .gnd(gnd), .vdd(vdd), .A(w_1_), .Y(_3458_) );
NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(e_reg_1_), .B(a_reg_28_), .Y(_3459_) );
INVX1 INVX1_484 ( .gnd(gnd), .vdd(vdd), .A(_3459_), .Y(_3460_) );
NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(e_reg_1_), .B(a_reg_28_), .Y(_3461_) );
NOR3X1 NOR3X1_60 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3461_), .C(_3460_), .Y(_3462_) );
INVX1 INVX1_485 ( .gnd(gnd), .vdd(vdd), .A(_3461_), .Y(_3463_) );
AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_3463_), .B(_3459_), .C(w_1_), .Y(_3464_) );
OAI21X1 OAI21X1_593 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_3464_), .C(_3457_), .Y(_3465_) );
INVX1 INVX1_486 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .Y(_3466_) );
NAND3X1 NAND3X1_85 ( .gnd(gnd), .vdd(vdd), .A(w_1_), .B(_3459_), .C(_3463_), .Y(_3467_) );
OAI21X1 OAI21X1_594 ( .gnd(gnd), .vdd(vdd), .A(_3461_), .B(_3460_), .C(_3458_), .Y(_3468_) );
NAND3X1 NAND3X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3467_), .B(_3468_), .C(_3466_), .Y(_3469_) );
NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_3469_), .B(_3465_), .Y(_3470_) );
NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3456_), .Y(_3471_) );
INVX4 INVX4_4 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf3), .Y(_3472_) );
NAND3X1 NAND3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3449_), .C(_3402_), .Y(_3473_) );
NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_3473_), .Y(_3474_) );
NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(d_reg_1_), .B(_3444_), .Y(_3475_) );
NAND3X1 NAND3X1_88 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_3438_), .C(_3441_), .Y(_3476_) );
NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_3476_), .B(_3475_), .Y(_3477_) );
OAI21X1 OAI21X1_595 ( .gnd(gnd), .vdd(vdd), .A(c_reg_1_), .B(b_reg_1_), .C(_3452_), .Y(_3478_) );
INVX1 INVX1_487 ( .gnd(gnd), .vdd(vdd), .A(_3454_), .Y(_3479_) );
OAI22X1 OAI22X1_43 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf2), .B(_3479_), .C(_3478_), .D(_3405__bF_buf3), .Y(_3480_) );
AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_3477_), .B(_3474__bF_buf4), .C(_3480_), .Y(_3481_) );
NAND3X1 NAND3X1_89 ( .gnd(gnd), .vdd(vdd), .A(_3457_), .B(_3468_), .C(_3467_), .Y(_3482_) );
OAI21X1 OAI21X1_596 ( .gnd(gnd), .vdd(vdd), .A(_3462_), .B(_3464_), .C(_3466_), .Y(_3483_) );
NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_3482_), .B(_3483_), .Y(_3484_) );
NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_3484_), .B(_3481_), .Y(_3485_) );
NAND3X1 NAND3X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_3485_), .C(_3425_), .Y(_3486_) );
NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_3470_), .B(_3481_), .Y(_3487_) );
NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_3484_), .B(_3456_), .Y(_3488_) );
NAND3X1 NAND3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3424_), .B(_3488_), .C(_3487_), .Y(_3489_) );
NAND3X1 NAND3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf2), .B(_3489_), .C(_3486_), .Y(_3490_) );
AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_3487_), .B(_3488_), .C(_3424_), .Y(_3491_) );
AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_3471_), .B(_3485_), .C(_3425_), .Y(_3492_) );
OAI21X1 OAI21X1_597 ( .gnd(gnd), .vdd(vdd), .A(_3491_), .B(_3492_), .C(_3472_), .Y(_3493_) );
NAND3X1 NAND3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .B(_3428_), .C(_3493_), .Y(_3494_) );
NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3427_), .Y(_3495_) );
NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_3490_), .B(_3493_), .Y(_3496_) );
AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_3496_), .B(_3495_), .C(_3385_), .Y(_3497_) );
INVX1 INVX1_488 ( .gnd(gnd), .vdd(vdd), .A(_3667__129_), .Y(_3498_) );
NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3432__bF_buf10), .Y(_3499_) );
AOI22X1 AOI22X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf10), .B(_3499_), .C(_3494_), .D(_3497_), .Y(_3500_) );
OAI21X1 OAI21X1_598 ( .gnd(gnd), .vdd(vdd), .A(_3436_), .B(_3387__bF_buf9), .C(_3500_), .Y(_5__1_) );
INVX1 INVX1_489 ( .gnd(gnd), .vdd(vdd), .A(a_reg_2_), .Y(_3501_) );
OAI21X1 OAI21X1_599 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_3492_), .C(_3486_), .Y(_3502_) );
OAI21X1 OAI21X1_600 ( .gnd(gnd), .vdd(vdd), .A(_3484_), .B(_3481_), .C(_3482_), .Y(_3503_) );
NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(c_reg_2_), .B(b_reg_2_), .Y(_3504_) );
NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(c_reg_2_), .B(b_reg_2_), .Y(_3505_) );
INVX1 INVX1_490 ( .gnd(gnd), .vdd(vdd), .A(_3505_), .Y(_3506_) );
NAND3X1 NAND3X1_94 ( .gnd(gnd), .vdd(vdd), .A(d_reg_2_), .B(_3504_), .C(_3506_), .Y(_3507_) );
INVX2 INVX2_9 ( .gnd(gnd), .vdd(vdd), .A(d_reg_2_), .Y(_3508_) );
INVX1 INVX1_491 ( .gnd(gnd), .vdd(vdd), .A(_3504_), .Y(_3509_) );
OAI21X1 OAI21X1_601 ( .gnd(gnd), .vdd(vdd), .A(_3505_), .B(_3509_), .C(_3508_), .Y(_3510_) );
AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_3507_), .B(_3510_), .Y(_3511_) );
AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3504_), .C(_3505_), .Y(_3512_) );
INVX1 INVX1_492 ( .gnd(gnd), .vdd(vdd), .A(_3512_), .Y(_3513_) );
OAI21X1 OAI21X1_602 ( .gnd(gnd), .vdd(vdd), .A(b_reg_2_), .B(_3508_), .C(_3504_), .Y(_3514_) );
INVX1 INVX1_493 ( .gnd(gnd), .vdd(vdd), .A(_3514_), .Y(_3515_) );
OAI22X1 OAI22X1_44 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf1), .B(_3515_), .C(_3405__bF_buf2), .D(_3513_), .Y(_3516_) );
AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_3511_), .B(_3474__bF_buf3), .C(_3516_), .Y(_3517_) );
OAI21X1 OAI21X1_603 ( .gnd(gnd), .vdd(vdd), .A(_3458_), .B(_3461_), .C(_3459_), .Y(_3518_) );
NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(e_reg_2_), .B(a_reg_29_), .Y(_3519_) );
NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(e_reg_2_), .B(a_reg_29_), .Y(_3520_) );
INVX1 INVX1_494 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .Y(_3521_) );
NAND3X1 NAND3X1_95 ( .gnd(gnd), .vdd(vdd), .A(w_2_), .B(_3519_), .C(_3521_), .Y(_3522_) );
INVX1 INVX1_495 ( .gnd(gnd), .vdd(vdd), .A(w_2_), .Y(_3523_) );
INVX1 INVX1_496 ( .gnd(gnd), .vdd(vdd), .A(_3519_), .Y(_3524_) );
OAI21X1 OAI21X1_604 ( .gnd(gnd), .vdd(vdd), .A(_3520_), .B(_3524_), .C(_3523_), .Y(_3525_) );
NAND3X1 NAND3X1_96 ( .gnd(gnd), .vdd(vdd), .A(_3518_), .B(_3525_), .C(_3522_), .Y(_3526_) );
INVX1 INVX1_497 ( .gnd(gnd), .vdd(vdd), .A(_3518_), .Y(_3527_) );
NOR3X1 NOR3X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3520_), .C(_3524_), .Y(_3528_) );
AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_3521_), .B(_3519_), .C(w_2_), .Y(_3529_) );
OAI21X1 OAI21X1_605 ( .gnd(gnd), .vdd(vdd), .A(_3528_), .B(_3529_), .C(_3527_), .Y(_3530_) );
NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3530_), .Y(_3531_) );
NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_3531_), .B(_3517_), .Y(_3532_) );
NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_3510_), .B(_3507_), .Y(_3533_) );
AOI22X1 AOI22X1_611 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf3), .B(_3514_), .C(_3451__bF_buf3), .D(_3512_), .Y(_3534_) );
OAI21X1 OAI21X1_606 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf2), .B(_3533_), .C(_3534_), .Y(_3535_) );
AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3530_), .C(_3535_), .Y(_3536_) );
OAI21X1 OAI21X1_607 ( .gnd(gnd), .vdd(vdd), .A(_3536_), .B(_3532_), .C(_3503_), .Y(_3537_) );
INVX1 INVX1_498 ( .gnd(gnd), .vdd(vdd), .A(_3482_), .Y(_3538_) );
AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_3456_), .B(_3470_), .C(_3538_), .Y(_3539_) );
NAND3X1 NAND3X1_97 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .B(_3530_), .C(_3535_), .Y(_3540_) );
NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_3531_), .B(_3517_), .Y(_3541_) );
NAND3X1 NAND3X1_98 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3541_), .C(_3539_), .Y(_3542_) );
AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_3542_), .B(_3537_), .C(_3392_), .Y(_3543_) );
NAND3X1 NAND3X1_99 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3541_), .C(_3503_), .Y(_3544_) );
OAI21X1 OAI21X1_608 ( .gnd(gnd), .vdd(vdd), .A(_3536_), .B(_3532_), .C(_3539_), .Y(_3545_) );
AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .B(_3545_), .C(_3391_), .Y(_3546_) );
OAI21X1 OAI21X1_609 ( .gnd(gnd), .vdd(vdd), .A(_3543_), .B(_3546_), .C(_3502_), .Y(_3547_) );
AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_3489_), .B(_3437__bF_buf1), .C(_3491_), .Y(_3548_) );
NAND3X1 NAND3X1_100 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .B(_3545_), .C(_3544_), .Y(_3549_) );
NAND3X1 NAND3X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3537_), .C(_3542_), .Y(_3550_) );
NAND3X1 NAND3X1_102 ( .gnd(gnd), .vdd(vdd), .A(_3548_), .B(_3549_), .C(_3550_), .Y(_3551_) );
AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3547_), .B(_3551_), .C(_3494_), .Y(_3552_) );
NAND3X1 NAND3X1_103 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_3489_), .C(_3486_), .Y(_3553_) );
OAI21X1 OAI21X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3491_), .B(_3492_), .C(_3437__bF_buf0), .Y(_3554_) );
AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_3554_), .B(_3553_), .C(_3495_), .Y(_3555_) );
NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_3551_), .B(_3547_), .Y(_3556_) );
OAI21X1 OAI21X1_611 ( .gnd(gnd), .vdd(vdd), .A(_3555_), .B(_3556_), .C(round_ctr_inc_bF_buf7), .Y(_3557_) );
NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3552_), .B(_3557_), .Y(_3558_) );
INVX1 INVX1_499 ( .gnd(gnd), .vdd(vdd), .A(_3667__130_), .Y(_3559_) );
NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .B(_3432__bF_buf9), .Y(_3560_) );
AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf9), .B(_3560_), .C(_3558_), .Y(_3561_) );
OAI21X1 OAI21X1_612 ( .gnd(gnd), .vdd(vdd), .A(_3501_), .B(_3387__bF_buf8), .C(_3561_), .Y(_5__2_) );
INVX1 INVX1_500 ( .gnd(gnd), .vdd(vdd), .A(a_reg_3_), .Y(_3562_) );
NAND3X1 NAND3X1_104 ( .gnd(gnd), .vdd(vdd), .A(_3549_), .B(_3550_), .C(_3502_), .Y(_3563_) );
OAI21X1 OAI21X1_613 ( .gnd(gnd), .vdd(vdd), .A(_3543_), .B(_3546_), .C(_3548_), .Y(_3564_) );
NAND3X1 NAND3X1_105 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .B(_3564_), .C(_3555_), .Y(_3565_) );
AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3540_), .B(_3541_), .C(_3503_), .Y(_3566_) );
OAI21X1 OAI21X1_614 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3566_), .C(_3544_), .Y(_3567_) );
OAI21X1 OAI21X1_615 ( .gnd(gnd), .vdd(vdd), .A(_3531_), .B(_3517_), .C(_3526_), .Y(_3568_) );
NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(c_reg_3_), .B(b_reg_3_), .Y(_3569_) );
INVX1 INVX1_501 ( .gnd(gnd), .vdd(vdd), .A(_3569_), .Y(_3570_) );
NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(c_reg_3_), .B(b_reg_3_), .Y(_3571_) );
OAI21X1 OAI21X1_616 ( .gnd(gnd), .vdd(vdd), .A(_3571_), .B(_3570_), .C(d_reg_3_), .Y(_3572_) );
INVX2 INVX2_10 ( .gnd(gnd), .vdd(vdd), .A(d_reg_3_), .Y(_3573_) );
INVX1 INVX1_502 ( .gnd(gnd), .vdd(vdd), .A(c_reg_3_), .Y(_3574_) );
INVX2 INVX2_11 ( .gnd(gnd), .vdd(vdd), .A(b_reg_3_), .Y(_3575_) );
NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_3575_), .Y(_3576_) );
NAND3X1 NAND3X1_106 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3569_), .C(_3576_), .Y(_3577_) );
AOI22X1 AOI22X1_612 ( .gnd(gnd), .vdd(vdd), .A(_3572_), .B(_3577_), .C(_3472_), .D(_3473_), .Y(_3578_) );
OAI21X1 OAI21X1_617 ( .gnd(gnd), .vdd(vdd), .A(d_reg_3_), .B(_3570_), .C(_3576_), .Y(_3579_) );
OAI21X1 OAI21X1_618 ( .gnd(gnd), .vdd(vdd), .A(b_reg_3_), .B(_3573_), .C(_3569_), .Y(_3580_) );
INVX1 INVX1_503 ( .gnd(gnd), .vdd(vdd), .A(_3580_), .Y(_3581_) );
OAI22X1 OAI22X1_45 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf0), .B(_3581_), .C(_3579_), .D(_3405__bF_buf1), .Y(_3582_) );
OAI21X1 OAI21X1_619 ( .gnd(gnd), .vdd(vdd), .A(_3523_), .B(_3520_), .C(_3519_), .Y(_3583_) );
INVX1 INVX1_504 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .Y(_3584_) );
NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(e_reg_3_), .B(a_reg_30_), .Y(_3585_) );
OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(e_reg_3_), .B(a_reg_30_), .Y(_3586_) );
NAND3X1 NAND3X1_107 ( .gnd(gnd), .vdd(vdd), .A(w_3_), .B(_3585_), .C(_3586_), .Y(_3587_) );
INVX1 INVX1_505 ( .gnd(gnd), .vdd(vdd), .A(w_3_), .Y(_3588_) );
INVX1 INVX1_506 ( .gnd(gnd), .vdd(vdd), .A(_3585_), .Y(_3589_) );
NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(e_reg_3_), .B(a_reg_30_), .Y(_3590_) );
OAI21X1 OAI21X1_620 ( .gnd(gnd), .vdd(vdd), .A(_3590_), .B(_3589_), .C(_3588_), .Y(_3591_) );
AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3587_), .B(_3591_), .C(_3584_), .Y(_3592_) );
NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_3587_), .B(_3591_), .Y(_3593_) );
NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .B(_3593_), .Y(_3594_) );
OAI22X1 OAI22X1_46 ( .gnd(gnd), .vdd(vdd), .A(_3578_), .B(_3582_), .C(_3592_), .D(_3594_), .Y(_3595_) );
NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_3577_), .B(_3572_), .Y(_3596_) );
AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf2), .B(_3596_), .C(_3582_), .Y(_3597_) );
NAND3X1 NAND3X1_108 ( .gnd(gnd), .vdd(vdd), .A(_3583_), .B(_3587_), .C(_3591_), .Y(_3598_) );
NOR3X1 NOR3X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(_3590_), .C(_3589_), .Y(_3599_) );
AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_3586_), .B(_3585_), .C(w_3_), .Y(_3600_) );
OAI21X1 OAI21X1_621 ( .gnd(gnd), .vdd(vdd), .A(_3600_), .B(_3599_), .C(_3584_), .Y(_3601_) );
NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .B(_3601_), .Y(_3602_) );
NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .B(_3597_), .Y(_3603_) );
NAND3X1 NAND3X1_109 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .B(_3603_), .C(_3568_), .Y(_3604_) );
INVX1 INVX1_507 ( .gnd(gnd), .vdd(vdd), .A(_3526_), .Y(_3605_) );
AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3535_), .B(_3530_), .C(_3605_), .Y(_3606_) );
NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .B(_3603_), .Y(_3607_) );
NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_3606_), .B(_3607_), .Y(_3608_) );
NAND3X1 NAND3X1_110 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf1), .B(_3604_), .C(_3608_), .Y(_3609_) );
OAI21X1 OAI21X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3605_), .B(_3532_), .C(_3607_), .Y(_3610_) );
NAND3X1 NAND3X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .B(_3603_), .C(_3606_), .Y(_3611_) );
NAND3X1 NAND3X1_112 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf1), .B(_3611_), .C(_3610_), .Y(_3612_) );
NAND3X1 NAND3X1_113 ( .gnd(gnd), .vdd(vdd), .A(_3609_), .B(_3612_), .C(_3567_), .Y(_3613_) );
INVX1 INVX1_508 ( .gnd(gnd), .vdd(vdd), .A(_3544_), .Y(_3614_) );
AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .B(_3545_), .C(_3614_), .Y(_3615_) );
AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_3610_), .B(_3611_), .C(_3474__bF_buf0), .Y(_3616_) );
AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3608_), .B(_3604_), .C(_3406__bF_buf0), .Y(_3617_) );
OAI21X1 OAI21X1_623 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3616_), .C(_3615_), .Y(_3618_) );
NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_3613_), .B(_3618_), .Y(_3619_) );
NAND3X1 NAND3X1_114 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .B(_3619_), .C(_3565_), .Y(_3620_) );
OAI21X1 OAI21X1_624 ( .gnd(gnd), .vdd(vdd), .A(_3617_), .B(_3616_), .C(_3567_), .Y(_3621_) );
NAND3X1 NAND3X1_115 ( .gnd(gnd), .vdd(vdd), .A(_3609_), .B(_3612_), .C(_3615_), .Y(_3622_) );
NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_3621_), .B(_3622_), .Y(_3623_) );
OAI21X1 OAI21X1_625 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .B(_3619_), .C(round_ctr_inc_bF_buf6), .Y(_3624_) );
AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3552_), .B(_3623_), .C(_3624_), .Y(_3625_) );
INVX1 INVX1_509 ( .gnd(gnd), .vdd(vdd), .A(_3667__131_), .Y(_3626_) );
NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_3432__bF_buf8), .Y(_3627_) );
AOI22X1 AOI22X1_613 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf8), .B(_3627_), .C(_3620_), .D(_3625_), .Y(_3628_) );
OAI21X1 OAI21X1_626 ( .gnd(gnd), .vdd(vdd), .A(_3562_), .B(_3387__bF_buf7), .C(_3628_), .Y(_5__3_) );
INVX1 INVX1_510 ( .gnd(gnd), .vdd(vdd), .A(a_reg_4_), .Y(_3629_) );
AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_3612_), .B(_3609_), .C(_3567_), .Y(_3630_) );
OAI21X1 OAI21X1_627 ( .gnd(gnd), .vdd(vdd), .A(_3563_), .B(_3630_), .C(_3613_), .Y(_3631_) );
AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_3552_), .B(_3623_), .C(_3631_), .Y(_3632_) );
NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3606_), .B(_3607_), .Y(_3633_) );
AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf4), .B(_3608_), .C(_3633_), .Y(_3634_) );
OAI21X1 OAI21X1_628 ( .gnd(gnd), .vdd(vdd), .A(_3602_), .B(_3597_), .C(_3598_), .Y(_3635_) );
AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(c_reg_4_), .B(b_reg_4_), .Y(_3636_) );
NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(c_reg_4_), .B(b_reg_4_), .Y(_3637_) );
OAI21X1 OAI21X1_629 ( .gnd(gnd), .vdd(vdd), .A(_3637_), .B(_3636_), .C(d_reg_4_), .Y(_3638_) );
INVX2 INVX2_12 ( .gnd(gnd), .vdd(vdd), .A(d_reg_4_), .Y(_3639_) );
NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(c_reg_4_), .B(b_reg_4_), .Y(_3640_) );
INVX1 INVX1_511 ( .gnd(gnd), .vdd(vdd), .A(c_reg_4_), .Y(_3641_) );
INVX1 INVX1_512 ( .gnd(gnd), .vdd(vdd), .A(b_reg_4_), .Y(_3642_) );
NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_3642_), .Y(_3643_) );
NAND3X1 NAND3X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(_3640_), .C(_3643_), .Y(_3644_) );
NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_3638_), .B(_3644_), .Y(_3645_) );
NAND3X1 NAND3X1_117 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf4), .B(_3405__bF_buf0), .C(_3645_), .Y(_3646_) );
AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(_3640_), .C(_3637_), .Y(_3647_) );
OAI21X1 OAI21X1_630 ( .gnd(gnd), .vdd(vdd), .A(b_reg_4_), .B(_3639_), .C(_3640_), .Y(_3648_) );
AOI22X1 AOI22X1_614 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf2), .B(_3648_), .C(_3451__bF_buf2), .D(_3647_), .Y(_3649_) );
OAI21X1 OAI21X1_631 ( .gnd(gnd), .vdd(vdd), .A(_3588_), .B(_3590_), .C(_3585_), .Y(_3650_) );
NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(e_reg_4_), .B(a_reg_31_), .Y(_3651_) );
OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(e_reg_4_), .B(a_reg_31_), .Y(_3652_) );
NAND3X1 NAND3X1_118 ( .gnd(gnd), .vdd(vdd), .A(w_4_), .B(_3651_), .C(_3652_), .Y(_3653_) );
INVX1 INVX1_513 ( .gnd(gnd), .vdd(vdd), .A(w_4_), .Y(_3654_) );
AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(e_reg_4_), .B(a_reg_31_), .Y(_3655_) );
NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(e_reg_4_), .B(a_reg_31_), .Y(_3656_) );
OAI21X1 OAI21X1_632 ( .gnd(gnd), .vdd(vdd), .A(_3656_), .B(_3655_), .C(_3654_), .Y(_3657_) );
NAND3X1 NAND3X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .B(_3657_), .C(_3653_), .Y(_3658_) );
INVX1 INVX1_514 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .Y(_3659_) );
NOR3X1 NOR3X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3654_), .B(_3656_), .C(_3655_), .Y(_3660_) );
AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_3652_), .B(_3651_), .C(w_4_), .Y(_3661_) );
OAI21X1 OAI21X1_633 ( .gnd(gnd), .vdd(vdd), .A(_3661_), .B(_3660_), .C(_3659_), .Y(_3662_) );
NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3662_), .Y(_3663_) );
AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_3646_), .B(_3649_), .C(_3663_), .Y(_3664_) );
AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_3644_), .B(_3638_), .Y(_12_) );
OAI21X1 OAI21X1_634 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf3), .B(_12_), .C(_3649_), .Y(_13_) );
AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .B(_3662_), .C(_13_), .Y(_14_) );
OAI21X1 OAI21X1_635 ( .gnd(gnd), .vdd(vdd), .A(_3664_), .B(_14_), .C(_3635_), .Y(_15_) );
AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_3572_), .B(_3577_), .Y(_16_) );
AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3569_), .C(_3571_), .Y(_17_) );
AOI22X1 AOI22X1_615 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf1), .B(_3580_), .C(_3451__bF_buf1), .D(_17_), .Y(_18_) );
OAI21X1 OAI21X1_636 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf2), .B(_16_), .C(_18_), .Y(_19_) );
INVX1 INVX1_515 ( .gnd(gnd), .vdd(vdd), .A(_3598_), .Y(_20_) );
AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_19_), .B(_3601_), .C(_20_), .Y(_21_) );
AOI22X1 AOI22X1_616 ( .gnd(gnd), .vdd(vdd), .A(_3638_), .B(_3644_), .C(_3472_), .D(_3473_), .Y(_22_) );
OAI21X1 OAI21X1_637 ( .gnd(gnd), .vdd(vdd), .A(d_reg_4_), .B(_3636_), .C(_3643_), .Y(_23_) );
INVX1 INVX1_516 ( .gnd(gnd), .vdd(vdd), .A(_3648_), .Y(_24_) );
OAI22X1 OAI22X1_47 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf3), .B(_24_), .C(_23_), .D(_3405__bF_buf5), .Y(_25_) );
AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_3653_), .B(_3657_), .C(_3659_), .Y(_26_) );
NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_3657_), .B(_3653_), .Y(_27_) );
NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(_3650_), .B(_27_), .Y(_28_) );
OAI22X1 OAI22X1_48 ( .gnd(gnd), .vdd(vdd), .A(_22_), .B(_25_), .C(_26_), .D(_28_), .Y(_29_) );
NAND3X1 NAND3X1_120 ( .gnd(gnd), .vdd(vdd), .A(_3646_), .B(_3649_), .C(_3663_), .Y(_30_) );
NAND3X1 NAND3X1_121 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .C(_21_), .Y(_31_) );
AOI22X1 AOI22X1_617 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3411__bF_buf2), .C(_15_), .D(_31_), .Y(_32_) );
NAND3X1 NAND3X1_122 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .C(_3635_), .Y(_33_) );
OAI21X1 OAI21X1_638 ( .gnd(gnd), .vdd(vdd), .A(_3664_), .B(_14_), .C(_21_), .Y(_34_) );
AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_33_), .B(_34_), .C(_3473_), .Y(_35_) );
OAI21X1 OAI21X1_639 ( .gnd(gnd), .vdd(vdd), .A(_32_), .B(_35_), .C(_3634_), .Y(_36_) );
AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_3595_), .B(_3603_), .C(_3568_), .Y(_37_) );
OAI21X1 OAI21X1_640 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf4), .B(_37_), .C(_3604_), .Y(_38_) );
NAND3X1 NAND3X1_123 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_34_), .C(_33_), .Y(_39_) );
INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .Y(_40_) );
NAND3X1 NAND3X1_124 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf3), .B(_15_), .C(_31_), .Y(_41_) );
NAND3X1 NAND3X1_125 ( .gnd(gnd), .vdd(vdd), .A(_39_), .B(_41_), .C(_38_), .Y(_42_) );
NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_42_), .B(_36_), .Y(_43_) );
OAI21X1 OAI21X1_641 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_3632_), .C(round_ctr_inc_bF_buf5), .Y(_44_) );
AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_3632_), .B(_43_), .C(_44_), .Y(_45_) );
INVX1 INVX1_517 ( .gnd(gnd), .vdd(vdd), .A(_3667__132_), .Y(_46_) );
NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_3432__bF_buf7), .Y(_47_) );
AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf7), .B(_47_), .C(_45_), .Y(_48_) );
OAI21X1 OAI21X1_642 ( .gnd(gnd), .vdd(vdd), .A(_3629_), .B(_3387__bF_buf6), .C(_48_), .Y(_5__4_) );
NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .Y(_49_) );
NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_49_), .Y(_50_) );
AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_34_), .C(_50_), .Y(_51_) );
AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf3), .B(_3645_), .C(_25_), .Y(_52_) );
OAI21X1 OAI21X1_643 ( .gnd(gnd), .vdd(vdd), .A(_3663_), .B(_52_), .C(_3658_), .Y(_53_) );
AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(c_reg_5_), .B(b_reg_5_), .Y(_54_) );
NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(c_reg_5_), .B(b_reg_5_), .Y(_55_) );
OAI21X1 OAI21X1_644 ( .gnd(gnd), .vdd(vdd), .A(_55_), .B(_54_), .C(d_reg_5_), .Y(_56_) );
INVX2 INVX2_13 ( .gnd(gnd), .vdd(vdd), .A(d_reg_5_), .Y(_57_) );
NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(c_reg_5_), .B(b_reg_5_), .Y(_58_) );
INVX1 INVX1_518 ( .gnd(gnd), .vdd(vdd), .A(c_reg_5_), .Y(_59_) );
INVX1 INVX1_519 ( .gnd(gnd), .vdd(vdd), .A(b_reg_5_), .Y(_60_) );
NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_60_), .Y(_61_) );
NAND3X1 NAND3X1_126 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .C(_61_), .Y(_62_) );
AOI22X1 AOI22X1_618 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_62_), .C(_3472_), .D(_3473_), .Y(_63_) );
AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_58_), .C(_55_), .Y(_64_) );
INVX1 INVX1_520 ( .gnd(gnd), .vdd(vdd), .A(_64_), .Y(_65_) );
OAI21X1 OAI21X1_645 ( .gnd(gnd), .vdd(vdd), .A(b_reg_5_), .B(_57_), .C(_58_), .Y(_66_) );
INVX1 INVX1_521 ( .gnd(gnd), .vdd(vdd), .A(_66_), .Y(_67_) );
OAI22X1 OAI22X1_49 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf1), .B(_67_), .C(_3405__bF_buf4), .D(_65_), .Y(_68_) );
OAI21X1 OAI21X1_646 ( .gnd(gnd), .vdd(vdd), .A(_3654_), .B(_3656_), .C(_3651_), .Y(_69_) );
INVX1 INVX1_522 ( .gnd(gnd), .vdd(vdd), .A(_69_), .Y(_70_) );
NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(a_reg_0_), .B(e_reg_5_), .Y(_71_) );
INVX2 INVX2_14 ( .gnd(gnd), .vdd(vdd), .A(e_reg_5_), .Y(_72_) );
NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_3384_), .B(_72_), .Y(_73_) );
NAND3X1 NAND3X1_127 ( .gnd(gnd), .vdd(vdd), .A(w_5_), .B(_71_), .C(_73_), .Y(_74_) );
INVX1 INVX1_523 ( .gnd(gnd), .vdd(vdd), .A(w_5_), .Y(_75_) );
AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(a_reg_0_), .B(e_reg_5_), .Y(_76_) );
NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(a_reg_0_), .B(e_reg_5_), .Y(_77_) );
OAI21X1 OAI21X1_647 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_76_), .C(_75_), .Y(_78_) );
AOI21X1 AOI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(_74_), .B(_78_), .C(_70_), .Y(_79_) );
NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_78_), .B(_74_), .Y(_80_) );
NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_80_), .Y(_81_) );
OAI22X1 OAI22X1_50 ( .gnd(gnd), .vdd(vdd), .A(_63_), .B(_68_), .C(_79_), .D(_81_), .Y(_82_) );
NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_56_), .B(_62_), .Y(_83_) );
NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_3474__bF_buf2), .Y(_84_) );
AOI22X1 AOI22X1_619 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf0), .B(_66_), .C(_3451__bF_buf0), .D(_64_), .Y(_85_) );
NAND3X1 NAND3X1_128 ( .gnd(gnd), .vdd(vdd), .A(_69_), .B(_78_), .C(_74_), .Y(_86_) );
NOR3X1 NOR3X1_64 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_77_), .C(_76_), .Y(_87_) );
AOI21X1 AOI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_71_), .C(w_5_), .Y(_88_) );
OAI21X1 OAI21X1_648 ( .gnd(gnd), .vdd(vdd), .A(_87_), .B(_88_), .C(_70_), .Y(_89_) );
NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_89_), .Y(_90_) );
NAND3X1 NAND3X1_129 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_84_), .C(_90_), .Y(_91_) );
NAND3X1 NAND3X1_130 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_91_), .C(_53_), .Y(_92_) );
INVX1 INVX1_524 ( .gnd(gnd), .vdd(vdd), .A(_3658_), .Y(_93_) );
AOI21X1 AOI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_13_), .B(_3662_), .C(_93_), .Y(_94_) );
AOI21X1 AOI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_84_), .B(_85_), .C(_90_), .Y(_95_) );
AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_62_), .B(_56_), .Y(_96_) );
OAI21X1 OAI21X1_649 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf1), .B(_96_), .C(_85_), .Y(_97_) );
AOI21X1 AOI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(_86_), .B(_89_), .C(_97_), .Y(_98_) );
OAI21X1 OAI21X1_650 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_98_), .C(_94_), .Y(_99_) );
AOI22X1 AOI22X1_620 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3411__bF_buf0), .C(_99_), .D(_92_), .Y(_100_) );
OAI21X1 OAI21X1_651 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_98_), .C(_53_), .Y(_101_) );
NAND3X1 NAND3X1_131 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_91_), .C(_94_), .Y(_102_) );
AOI21X1 AOI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_101_), .C(_3473_), .Y(_103_) );
OAI21X1 OAI21X1_652 ( .gnd(gnd), .vdd(vdd), .A(_100_), .B(_103_), .C(_51_), .Y(_104_) );
AOI21X1 AOI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_29_), .B(_30_), .C(_3635_), .Y(_105_) );
OAI21X1 OAI21X1_653 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf2), .B(_105_), .C(_33_), .Y(_106_) );
NAND3X1 NAND3X1_132 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_101_), .C(_102_), .Y(_107_) );
NAND3X1 NAND3X1_133 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf1), .B(_99_), .C(_92_), .Y(_108_) );
NAND3X1 NAND3X1_134 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_108_), .C(_106_), .Y(_109_) );
NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_104_), .Y(_110_) );
OAI21X1 OAI21X1_654 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_3632_), .C(_42_), .Y(_111_) );
XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_111_), .B(_110_), .Y(_112_) );
INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(_3387__bF_buf5), .Y(_113_) );
INVX1 INVX1_525 ( .gnd(gnd), .vdd(vdd), .A(_3667__133_), .Y(_114_) );
NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_3432__bF_buf6), .Y(_115_) );
AOI22X1 AOI22X1_621 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_3433__bF_buf6), .C(a_reg_5_), .D(_113__bF_buf4), .Y(_116_) );
OAI21X1 OAI21X1_655 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_112_), .C(_116_), .Y(_5__5_) );
NOR3X1 NOR3X1_65 ( .gnd(gnd), .vdd(vdd), .A(_3548_), .B(_3543_), .C(_3546_), .Y(_117_) );
INVX1 INVX1_526 ( .gnd(gnd), .vdd(vdd), .A(_3613_), .Y(_118_) );
AOI21X1 AOI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_3618_), .C(_118_), .Y(_119_) );
OAI21X1 OAI21X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3565_), .B(_3619_), .C(_119_), .Y(_120_) );
NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_43_), .Y(_121_) );
NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_120_), .Y(_122_) );
AOI21X1 AOI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_108_), .C(_106_), .Y(_123_) );
OAI21X1 OAI21X1_657 ( .gnd(gnd), .vdd(vdd), .A(_123_), .B(_42_), .C(_109_), .Y(_124_) );
INVX1 INVX1_527 ( .gnd(gnd), .vdd(vdd), .A(_124_), .Y(_125_) );
NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_91_), .Y(_126_) );
NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_126_), .Y(_127_) );
AOI21X1 AOI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf0), .B(_99_), .C(_127_), .Y(_128_) );
AOI21X1 AOI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf1), .B(_83_), .C(_68_), .Y(_129_) );
OAI21X1 OAI21X1_658 ( .gnd(gnd), .vdd(vdd), .A(_90_), .B(_129_), .C(_86_), .Y(_130_) );
INVX2 INVX2_15 ( .gnd(gnd), .vdd(vdd), .A(d_reg_6_), .Y(_131_) );
NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(c_reg_6_), .B(b_reg_6_), .Y(_132_) );
NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_132_), .Y(_133_) );
NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(c_reg_6_), .B(b_reg_6_), .Y(_134_) );
AOI21X1 AOI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_134_), .C(_132_), .Y(_135_) );
OAI21X1 OAI21X1_659 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_134_), .C(_135_), .Y(_136_) );
NAND3X1 NAND3X1_135 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_136_), .C(_3474__bF_buf0), .Y(_137_) );
OAI21X1 OAI21X1_660 ( .gnd(gnd), .vdd(vdd), .A(b_reg_6_), .B(_131_), .C(_134_), .Y(_138_) );
AOI22X1 AOI22X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf4), .B(_138_), .C(_3451__bF_buf4), .D(_135_), .Y(_139_) );
OAI21X1 OAI21X1_661 ( .gnd(gnd), .vdd(vdd), .A(_75_), .B(_77_), .C(_71_), .Y(_140_) );
INVX1 INVX1_528 ( .gnd(gnd), .vdd(vdd), .A(w_6_), .Y(_141_) );
NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(a_reg_1_), .B(e_reg_6_), .Y(_142_) );
INVX1 INVX1_529 ( .gnd(gnd), .vdd(vdd), .A(_142_), .Y(_143_) );
NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(a_reg_1_), .B(e_reg_6_), .Y(_144_) );
NOR3X1 NOR3X1_66 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_144_), .C(_143_), .Y(_145_) );
INVX1 INVX1_530 ( .gnd(gnd), .vdd(vdd), .A(_144_), .Y(_146_) );
AOI21X1 AOI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(_146_), .B(_142_), .C(w_6_), .Y(_147_) );
OAI21X1 OAI21X1_662 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_147_), .C(_140_), .Y(_148_) );
INVX1 INVX1_531 ( .gnd(gnd), .vdd(vdd), .A(_140_), .Y(_149_) );
NAND3X1 NAND3X1_136 ( .gnd(gnd), .vdd(vdd), .A(w_6_), .B(_142_), .C(_146_), .Y(_150_) );
OAI21X1 OAI21X1_663 ( .gnd(gnd), .vdd(vdd), .A(_144_), .B(_143_), .C(_141_), .Y(_151_) );
NAND3X1 NAND3X1_137 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_151_), .C(_149_), .Y(_152_) );
AOI22X1 AOI22X1_623 ( .gnd(gnd), .vdd(vdd), .A(_148_), .B(_152_), .C(_139_), .D(_137_), .Y(_153_) );
NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_136_), .Y(_154_) );
OAI21X1 OAI21X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf0), .B(_154_), .C(_139_), .Y(_155_) );
NAND3X1 NAND3X1_138 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_151_), .C(_150_), .Y(_156_) );
OAI21X1 OAI21X1_665 ( .gnd(gnd), .vdd(vdd), .A(_145_), .B(_147_), .C(_149_), .Y(_157_) );
AOI21X1 AOI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .C(_155_), .Y(_158_) );
OAI21X1 OAI21X1_666 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_158_), .C(_130_), .Y(_159_) );
INVX1 INVX1_532 ( .gnd(gnd), .vdd(vdd), .A(_86_), .Y(_160_) );
AOI21X1 AOI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_89_), .C(_160_), .Y(_161_) );
NAND3X1 NAND3X1_139 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .C(_155_), .Y(_162_) );
NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_157_), .Y(_163_) );
NAND3X1 NAND3X1_140 ( .gnd(gnd), .vdd(vdd), .A(_137_), .B(_139_), .C(_163_), .Y(_164_) );
NAND3X1 NAND3X1_141 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_164_), .C(_161_), .Y(_165_) );
AOI22X1 AOI22X1_624 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3449_), .C(_165_), .D(_159_), .Y(_166_) );
NAND3X1 NAND3X1_142 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_164_), .C(_130_), .Y(_167_) );
OAI21X1 OAI21X1_667 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_158_), .C(_161_), .Y(_168_) );
AOI21X1 AOI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_168_), .C(_3391_), .Y(_169_) );
OAI21X1 OAI21X1_668 ( .gnd(gnd), .vdd(vdd), .A(_166_), .B(_169_), .C(_128_), .Y(_170_) );
AOI21X1 AOI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(_82_), .B(_91_), .C(_53_), .Y(_171_) );
OAI21X1 OAI21X1_669 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_171_), .C(_92_), .Y(_172_) );
NAND3X1 NAND3X1_143 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .B(_168_), .C(_167_), .Y(_173_) );
NAND3X1 NAND3X1_144 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_165_), .C(_159_), .Y(_174_) );
NAND3X1 NAND3X1_145 ( .gnd(gnd), .vdd(vdd), .A(_174_), .B(_173_), .C(_172_), .Y(_175_) );
NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_170_), .Y(_176_) );
AOI21X1 AOI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_122_), .B(_125_), .C(_176_), .Y(_177_) );
NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_125_), .B(_122_), .Y(_178_) );
INVX1 INVX1_533 ( .gnd(gnd), .vdd(vdd), .A(_176_), .Y(_179_) );
OAI21X1 OAI21X1_670 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_178_), .C(round_ctr_inc_bF_buf4), .Y(_180_) );
INVX1 INVX1_534 ( .gnd(gnd), .vdd(vdd), .A(_3667__134_), .Y(_181_) );
NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_3432__bF_buf5), .Y(_182_) );
AOI22X1 AOI22X1_625 ( .gnd(gnd), .vdd(vdd), .A(_182_), .B(_3433__bF_buf5), .C(a_reg_6_), .D(_113__bF_buf3), .Y(_183_) );
OAI21X1 OAI21X1_671 ( .gnd(gnd), .vdd(vdd), .A(_177_), .B(_180_), .C(_183_), .Y(_5__6_) );
INVX1 INVX1_535 ( .gnd(gnd), .vdd(vdd), .A(_175_), .Y(_184_) );
NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_184_), .B(_177_), .Y(_185_) );
NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_173_), .Y(_186_) );
NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_156_), .B(_162_), .Y(_187_) );
NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(c_reg_7_), .B(b_reg_7_), .Y(_188_) );
INVX2 INVX2_16 ( .gnd(gnd), .vdd(vdd), .A(c_reg_7_), .Y(_189_) );
INVX1 INVX1_536 ( .gnd(gnd), .vdd(vdd), .A(b_reg_7_), .Y(_190_) );
NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_190_), .Y(_191_) );
NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_191_), .Y(_192_) );
NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(d_reg_7_), .B(_192_), .Y(_193_) );
INVX2 INVX2_17 ( .gnd(gnd), .vdd(vdd), .A(d_reg_7_), .Y(_194_) );
NAND3X1 NAND3X1_146 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_188_), .C(_191_), .Y(_195_) );
NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_193_), .Y(_196_) );
OAI21X1 OAI21X1_672 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_190_), .C(_194_), .Y(_197_) );
OAI21X1 OAI21X1_673 ( .gnd(gnd), .vdd(vdd), .A(c_reg_7_), .B(b_reg_7_), .C(_197_), .Y(_198_) );
NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(b_reg_7_), .B(_189_), .Y(_199_) );
OAI21X1 OAI21X1_674 ( .gnd(gnd), .vdd(vdd), .A(b_reg_7_), .B(d_reg_7_), .C(_199_), .Y(_200_) );
OAI22X1 OAI22X1_51 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf4), .B(_200_), .C(_198_), .D(_3405__bF_buf3), .Y(_201_) );
AOI21X1 AOI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_196_), .B(_3474__bF_buf4), .C(_201_), .Y(_202_) );
OAI21X1 OAI21X1_675 ( .gnd(gnd), .vdd(vdd), .A(_141_), .B(_144_), .C(_142_), .Y(_203_) );
INVX2 INVX2_18 ( .gnd(gnd), .vdd(vdd), .A(w_7_), .Y(_204_) );
NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(a_reg_2_), .B(e_reg_7_), .Y(_205_) );
INVX1 INVX1_537 ( .gnd(gnd), .vdd(vdd), .A(e_reg_7_), .Y(_206_) );
NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_3501_), .B(_206_), .Y(_207_) );
NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_207_), .Y(_208_) );
OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_208_), .B(_204_), .Y(_209_) );
INVX1 INVX1_538 ( .gnd(gnd), .vdd(vdd), .A(_205_), .Y(_210_) );
NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(a_reg_2_), .B(e_reg_7_), .Y(_211_) );
OAI21X1 OAI21X1_676 ( .gnd(gnd), .vdd(vdd), .A(_211_), .B(_210_), .C(_204_), .Y(_212_) );
NAND3X1 NAND3X1_147 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_212_), .C(_209_), .Y(_213_) );
INVX1 INVX1_539 ( .gnd(gnd), .vdd(vdd), .A(_203_), .Y(_214_) );
NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_208_), .Y(_215_) );
INVX1 INVX1_540 ( .gnd(gnd), .vdd(vdd), .A(_212_), .Y(_216_) );
OAI21X1 OAI21X1_677 ( .gnd(gnd), .vdd(vdd), .A(_215_), .B(_216_), .C(_214_), .Y(_217_) );
NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_217_), .B(_213_), .Y(_218_) );
NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_218_), .Y(_219_) );
INVX1 INVX1_541 ( .gnd(gnd), .vdd(vdd), .A(_219_), .Y(_220_) );
NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_218_), .Y(_221_) );
NAND3X1 NAND3X1_148 ( .gnd(gnd), .vdd(vdd), .A(_221_), .B(_187_), .C(_220_), .Y(_222_) );
INVX1 INVX1_542 ( .gnd(gnd), .vdd(vdd), .A(_187_), .Y(_223_) );
INVX1 INVX1_543 ( .gnd(gnd), .vdd(vdd), .A(_221_), .Y(_224_) );
OAI21X1 OAI21X1_678 ( .gnd(gnd), .vdd(vdd), .A(_219_), .B(_224_), .C(_223_), .Y(_225_) );
NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_225_), .Y(_226_) );
NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_186_), .B(_226_), .Y(_227_) );
OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_226_), .B(_186_), .Y(_228_) );
NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_227_), .B(_228_), .Y(_229_) );
AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_229_), .Y(_230_) );
OAI21X1 OAI21X1_679 ( .gnd(gnd), .vdd(vdd), .A(_229_), .B(_185_), .C(round_ctr_inc_bF_buf3), .Y(_231_) );
INVX1 INVX1_544 ( .gnd(gnd), .vdd(vdd), .A(_3667__135_), .Y(_232_) );
NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_3432__bF_buf4), .Y(_233_) );
AOI22X1 AOI22X1_626 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_3433__bF_buf4), .C(a_reg_7_), .D(_113__bF_buf2), .Y(_234_) );
OAI21X1 OAI21X1_680 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .C(_234_), .Y(_5__7_) );
NAND3X1 NAND3X1_149 ( .gnd(gnd), .vdd(vdd), .A(_222_), .B(_225_), .C(_186_), .Y(_235_) );
NAND3X1 NAND3X1_150 ( .gnd(gnd), .vdd(vdd), .A(_167_), .B(_173_), .C(_226_), .Y(_236_) );
AOI21X1 AOI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_235_), .B(_236_), .C(_176_), .Y(_237_) );
NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(_237_), .B(_121_), .Y(_238_) );
NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_175_), .B(_227_), .Y(_239_) );
AOI22X1 AOI22X1_627 ( .gnd(gnd), .vdd(vdd), .A(_228_), .B(_239_), .C(_124_), .D(_237_), .Y(_240_) );
OAI21X1 OAI21X1_681 ( .gnd(gnd), .vdd(vdd), .A(_3632_), .B(_238_), .C(_240_), .Y(_241_) );
INVX2 INVX2_19 ( .gnd(gnd), .vdd(vdd), .A(_241_), .Y(_242_) );
INVX1 INVX1_545 ( .gnd(gnd), .vdd(vdd), .A(_213_), .Y(_243_) );
NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(c_reg_8_), .B(b_reg_8_), .Y(_244_) );
INVX1 INVX1_546 ( .gnd(gnd), .vdd(vdd), .A(_244_), .Y(_245_) );
NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(c_reg_8_), .B(b_reg_8_), .Y(_246_) );
OAI21X1 OAI21X1_682 ( .gnd(gnd), .vdd(vdd), .A(_246_), .B(_245_), .C(d_reg_8_), .Y(_247_) );
INVX2 INVX2_20 ( .gnd(gnd), .vdd(vdd), .A(d_reg_8_), .Y(_248_) );
INVX1 INVX1_547 ( .gnd(gnd), .vdd(vdd), .A(_246_), .Y(_249_) );
NAND3X1 NAND3X1_151 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_244_), .C(_249_), .Y(_250_) );
AOI21X1 AOI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_250_), .C(_3406__bF_buf4), .Y(_251_) );
AOI21X1 AOI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_244_), .C(_246_), .Y(_252_) );
NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_3451__bF_buf3), .Y(_253_) );
INVX1 INVX1_548 ( .gnd(gnd), .vdd(vdd), .A(c_reg_8_), .Y(_254_) );
NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(b_reg_8_), .B(_254_), .Y(_255_) );
OAI21X1 OAI21X1_683 ( .gnd(gnd), .vdd(vdd), .A(b_reg_8_), .B(d_reg_8_), .C(_255_), .Y(_256_) );
OAI21X1 OAI21X1_684 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf3), .B(_256_), .C(_253_), .Y(_257_) );
OAI21X1 OAI21X1_685 ( .gnd(gnd), .vdd(vdd), .A(_204_), .B(_211_), .C(_205_), .Y(_258_) );
NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(a_reg_3_), .B(e_reg_8_), .Y(_259_) );
NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(a_reg_3_), .B(e_reg_8_), .Y(_260_) );
INVX1 INVX1_549 ( .gnd(gnd), .vdd(vdd), .A(_260_), .Y(_261_) );
NAND3X1 NAND3X1_152 ( .gnd(gnd), .vdd(vdd), .A(w_8_), .B(_259_), .C(_261_), .Y(_262_) );
INVX1 INVX1_550 ( .gnd(gnd), .vdd(vdd), .A(w_8_), .Y(_263_) );
INVX1 INVX1_551 ( .gnd(gnd), .vdd(vdd), .A(_259_), .Y(_264_) );
OAI21X1 OAI21X1_686 ( .gnd(gnd), .vdd(vdd), .A(_260_), .B(_264_), .C(_263_), .Y(_265_) );
NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(_265_), .B(_262_), .Y(_266_) );
NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_266_), .Y(_267_) );
INVX1 INVX1_552 ( .gnd(gnd), .vdd(vdd), .A(_258_), .Y(_268_) );
AOI21X1 AOI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_262_), .B(_265_), .C(_268_), .Y(_269_) );
OAI22X1 OAI22X1_52 ( .gnd(gnd), .vdd(vdd), .A(_267_), .B(_269_), .C(_257_), .D(_251_), .Y(_270_) );
NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_247_), .B(_250_), .Y(_271_) );
OAI21X1 OAI21X1_687 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf3), .B(_40__bF_buf3), .C(_271_), .Y(_272_) );
NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf2), .B(_256_), .Y(_273_) );
AOI21X1 AOI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf2), .B(_252_), .C(_273_), .Y(_274_) );
NAND3X1 NAND3X1_153 ( .gnd(gnd), .vdd(vdd), .A(_258_), .B(_265_), .C(_262_), .Y(_275_) );
NOR3X1 NOR3X1_67 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_260_), .C(_264_), .Y(_276_) );
AOI21X1 AOI21X1_73 ( .gnd(gnd), .vdd(vdd), .A(_261_), .B(_259_), .C(w_8_), .Y(_277_) );
OAI21X1 OAI21X1_688 ( .gnd(gnd), .vdd(vdd), .A(_276_), .B(_277_), .C(_268_), .Y(_278_) );
NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_278_), .Y(_279_) );
NAND3X1 NAND3X1_154 ( .gnd(gnd), .vdd(vdd), .A(_274_), .B(_272_), .C(_279_), .Y(_280_) );
NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_280_), .Y(_281_) );
OAI21X1 OAI21X1_689 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_219_), .C(_281_), .Y(_282_) );
AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_193_), .B(_195_), .Y(_283_) );
INVX1 INVX1_553 ( .gnd(gnd), .vdd(vdd), .A(_201_), .Y(_284_) );
OAI21X1 OAI21X1_690 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf3), .B(_283_), .C(_284_), .Y(_285_) );
AOI21X1 AOI21X1_74 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_217_), .C(_243_), .Y(_286_) );
NAND3X1 NAND3X1_155 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_280_), .C(_286_), .Y(_287_) );
AOI21X1 AOI21X1_75 ( .gnd(gnd), .vdd(vdd), .A(_287_), .B(_282_), .C(_3451__bF_buf1), .Y(_288_) );
OAI21X1 OAI21X1_691 ( .gnd(gnd), .vdd(vdd), .A(_202_), .B(_218_), .C(_213_), .Y(_289_) );
NAND3X1 NAND3X1_156 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_280_), .C(_289_), .Y(_290_) );
NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_286_), .Y(_291_) );
AOI21X1 AOI21X1_76 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_290_), .C(_3405__bF_buf2), .Y(_292_) );
OAI21X1 OAI21X1_692 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_288_), .C(_225_), .Y(_293_) );
AOI21X1 AOI21X1_77 ( .gnd(gnd), .vdd(vdd), .A(_220_), .B(_221_), .C(_187_), .Y(_294_) );
NAND3X1 NAND3X1_157 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf1), .B(_290_), .C(_291_), .Y(_295_) );
NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_281_), .B(_286_), .Y(_296_) );
AOI21X1 AOI21X1_78 ( .gnd(gnd), .vdd(vdd), .A(_270_), .B(_280_), .C(_289_), .Y(_297_) );
OAI21X1 OAI21X1_693 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_296_), .C(_3451__bF_buf0), .Y(_298_) );
NAND3X1 NAND3X1_158 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_295_), .C(_298_), .Y(_299_) );
AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_299_), .Y(_300_) );
OAI21X1 OAI21X1_694 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_242_), .C(round_ctr_inc_bF_buf2), .Y(_301_) );
AOI21X1 AOI21X1_79 ( .gnd(gnd), .vdd(vdd), .A(_242_), .B(_300_), .C(_301_), .Y(_302_) );
INVX1 INVX1_554 ( .gnd(gnd), .vdd(vdd), .A(a_reg_8_), .Y(_303_) );
OAI21X1 OAI21X1_695 ( .gnd(gnd), .vdd(vdd), .A(_3667__136_), .B(_3432__bF_buf3), .C(_3433__bF_buf3), .Y(_304_) );
OAI21X1 OAI21X1_696 ( .gnd(gnd), .vdd(vdd), .A(_303_), .B(_3387__bF_buf4), .C(_304_), .Y(_305_) );
OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_302_), .B(_305_), .Y(_5__8_) );
INVX1 INVX1_555 ( .gnd(gnd), .vdd(vdd), .A(a_reg_9_), .Y(_306_) );
OAI21X1 OAI21X1_697 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf4), .B(_297_), .C(_290_), .Y(_307_) );
AOI21X1 AOI21X1_80 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf3), .B(_271_), .C(_257_), .Y(_308_) );
OAI21X1 OAI21X1_698 ( .gnd(gnd), .vdd(vdd), .A(_279_), .B(_308_), .C(_275_), .Y(_309_) );
INVX2 INVX2_21 ( .gnd(gnd), .vdd(vdd), .A(d_reg_9_), .Y(_310_) );
NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(c_reg_9_), .B(b_reg_9_), .Y(_311_) );
INVX2 INVX2_22 ( .gnd(gnd), .vdd(vdd), .A(c_reg_9_), .Y(_312_) );
INVX2 INVX2_23 ( .gnd(gnd), .vdd(vdd), .A(b_reg_9_), .Y(_313_) );
NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_313_), .Y(_314_) );
NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(_311_), .B(_314_), .Y(_315_) );
XNOR2X1 XNOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(_310_), .Y(_316_) );
OAI21X1 OAI21X1_699 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_313_), .C(_310_), .Y(_317_) );
AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_317_), .B(_314_), .Y(_318_) );
NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(b_reg_9_), .B(_312_), .Y(_319_) );
OAI21X1 OAI21X1_700 ( .gnd(gnd), .vdd(vdd), .A(b_reg_9_), .B(d_reg_9_), .C(_319_), .Y(_320_) );
NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf1), .B(_320_), .Y(_321_) );
AOI21X1 AOI21X1_81 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf3), .B(_318_), .C(_321_), .Y(_322_) );
OAI21X1 OAI21X1_701 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf2), .B(_316_), .C(_322_), .Y(_323_) );
OAI21X1 OAI21X1_702 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_260_), .C(_259_), .Y(_324_) );
NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(a_reg_4_), .B(e_reg_9_), .Y(_325_) );
NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(a_reg_4_), .B(e_reg_9_), .Y(_326_) );
INVX1 INVX1_556 ( .gnd(gnd), .vdd(vdd), .A(_326_), .Y(_327_) );
NAND3X1 NAND3X1_159 ( .gnd(gnd), .vdd(vdd), .A(w_9_), .B(_325_), .C(_327_), .Y(_328_) );
INVX1 INVX1_557 ( .gnd(gnd), .vdd(vdd), .A(w_9_), .Y(_329_) );
INVX1 INVX1_558 ( .gnd(gnd), .vdd(vdd), .A(_325_), .Y(_330_) );
OAI21X1 OAI21X1_703 ( .gnd(gnd), .vdd(vdd), .A(_326_), .B(_330_), .C(_329_), .Y(_331_) );
NAND3X1 NAND3X1_160 ( .gnd(gnd), .vdd(vdd), .A(_324_), .B(_331_), .C(_328_), .Y(_332_) );
INVX1 INVX1_559 ( .gnd(gnd), .vdd(vdd), .A(_324_), .Y(_333_) );
NOR3X1 NOR3X1_68 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_326_), .C(_330_), .Y(_334_) );
AOI21X1 AOI21X1_82 ( .gnd(gnd), .vdd(vdd), .A(_327_), .B(_325_), .C(w_9_), .Y(_335_) );
OAI21X1 OAI21X1_704 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_335_), .C(_333_), .Y(_336_) );
AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_336_), .B(_332_), .Y(_337_) );
NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_323_), .Y(_338_) );
XNOR2X1 XNOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_315_), .B(d_reg_9_), .Y(_339_) );
OAI21X1 OAI21X1_705 ( .gnd(gnd), .vdd(vdd), .A(c_reg_9_), .B(b_reg_9_), .C(_317_), .Y(_340_) );
OAI22X1 OAI22X1_53 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf0), .B(_320_), .C(_340_), .D(_3405__bF_buf0), .Y(_341_) );
AOI21X1 AOI21X1_83 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_3474__bF_buf2), .C(_341_), .Y(_342_) );
NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_332_), .B(_336_), .Y(_343_) );
NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_342_), .Y(_344_) );
NAND3X1 NAND3X1_161 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_344_), .C(_309_), .Y(_345_) );
INVX1 INVX1_560 ( .gnd(gnd), .vdd(vdd), .A(_271_), .Y(_346_) );
OAI21X1 OAI21X1_706 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf1), .B(_346_), .C(_274_), .Y(_347_) );
INVX1 INVX1_561 ( .gnd(gnd), .vdd(vdd), .A(_275_), .Y(_348_) );
AOI21X1 AOI21X1_84 ( .gnd(gnd), .vdd(vdd), .A(_347_), .B(_278_), .C(_348_), .Y(_349_) );
NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_342_), .Y(_350_) );
NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_337_), .B(_323_), .Y(_351_) );
OAI21X1 OAI21X1_707 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_350_), .C(_349_), .Y(_352_) );
AOI22X1 AOI22X1_628 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3411__bF_buf4), .C(_352_), .D(_345_), .Y(_353_) );
OAI21X1 OAI21X1_708 ( .gnd(gnd), .vdd(vdd), .A(_351_), .B(_350_), .C(_309_), .Y(_354_) );
NAND3X1 NAND3X1_162 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_344_), .C(_349_), .Y(_355_) );
AOI21X1 AOI21X1_85 ( .gnd(gnd), .vdd(vdd), .A(_354_), .B(_355_), .C(_3473_), .Y(_356_) );
OAI21X1 OAI21X1_709 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_356_), .C(_307_), .Y(_357_) );
AOI21X1 AOI21X1_86 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf5), .B(_291_), .C(_296_), .Y(_358_) );
NAND3X1 NAND3X1_163 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_355_), .C(_354_), .Y(_359_) );
NAND3X1 NAND3X1_164 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf2), .B(_352_), .C(_345_), .Y(_360_) );
NAND3X1 NAND3X1_165 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_360_), .C(_358_), .Y(_361_) );
NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_361_), .B(_357_), .Y(_362_) );
NAND3X1 NAND3X1_166 ( .gnd(gnd), .vdd(vdd), .A(_225_), .B(_295_), .C(_298_), .Y(_363_) );
OAI21X1 OAI21X1_710 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_242_), .C(_363_), .Y(_364_) );
XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_364_), .B(_362_), .Y(_365_) );
INVX1 INVX1_562 ( .gnd(gnd), .vdd(vdd), .A(_3667__137_), .Y(_366_) );
OAI21X1 OAI21X1_711 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_366_), .Y(_367_) );
AOI22X1 AOI22X1_629 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf2), .B(_367_), .C(round_ctr_inc_bF_buf1), .D(_365_), .Y(_368_) );
OAI21X1 OAI21X1_712 ( .gnd(gnd), .vdd(vdd), .A(_306_), .B(_3387__bF_buf3), .C(_368_), .Y(_5__9_) );
AOI22X1 AOI22X1_630 ( .gnd(gnd), .vdd(vdd), .A(_357_), .B(_361_), .C(_299_), .D(_293_), .Y(_369_) );
NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_241_), .Y(_370_) );
NAND3X1 NAND3X1_167 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_360_), .C(_307_), .Y(_371_) );
AOI21X1 AOI21X1_87 ( .gnd(gnd), .vdd(vdd), .A(_360_), .B(_359_), .C(_307_), .Y(_372_) );
OAI21X1 OAI21X1_713 ( .gnd(gnd), .vdd(vdd), .A(_372_), .B(_363_), .C(_371_), .Y(_373_) );
INVX1 INVX1_563 ( .gnd(gnd), .vdd(vdd), .A(_373_), .Y(_374_) );
NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_370_), .Y(_375_) );
AOI21X1 AOI21X1_88 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_344_), .C(_309_), .Y(_376_) );
OAI21X1 OAI21X1_714 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_376_), .C(_345_), .Y(_377_) );
INVX1 INVX1_564 ( .gnd(gnd), .vdd(vdd), .A(_332_), .Y(_378_) );
NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(c_reg_10_), .B(b_reg_10_), .Y(_379_) );
INVX1 INVX1_565 ( .gnd(gnd), .vdd(vdd), .A(_379_), .Y(_380_) );
NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(c_reg_10_), .B(b_reg_10_), .Y(_381_) );
OAI21X1 OAI21X1_715 ( .gnd(gnd), .vdd(vdd), .A(_381_), .B(_380_), .C(d_reg_10_), .Y(_382_) );
INVX2 INVX2_24 ( .gnd(gnd), .vdd(vdd), .A(d_reg_10_), .Y(_383_) );
INVX1 INVX1_566 ( .gnd(gnd), .vdd(vdd), .A(_381_), .Y(_384_) );
NAND3X1 NAND3X1_168 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_379_), .C(_384_), .Y(_385_) );
AOI21X1 AOI21X1_89 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_385_), .C(_3406__bF_buf0), .Y(_386_) );
AOI21X1 AOI21X1_90 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_379_), .C(_381_), .Y(_387_) );
NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_3451__bF_buf2), .Y(_388_) );
INVX2 INVX2_25 ( .gnd(gnd), .vdd(vdd), .A(c_reg_10_), .Y(_389_) );
NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(b_reg_10_), .B(_389_), .Y(_390_) );
OAI21X1 OAI21X1_716 ( .gnd(gnd), .vdd(vdd), .A(b_reg_10_), .B(d_reg_10_), .C(_390_), .Y(_391_) );
OAI21X1 OAI21X1_717 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf3), .B(_391_), .C(_388_), .Y(_392_) );
OAI21X1 OAI21X1_718 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_326_), .C(_325_), .Y(_393_) );
INVX1 INVX1_567 ( .gnd(gnd), .vdd(vdd), .A(_393_), .Y(_394_) );
NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(a_reg_5_), .B(e_reg_10_), .Y(_395_) );
NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(a_reg_5_), .B(e_reg_10_), .Y(_396_) );
INVX1 INVX1_568 ( .gnd(gnd), .vdd(vdd), .A(_396_), .Y(_397_) );
NAND3X1 NAND3X1_169 ( .gnd(gnd), .vdd(vdd), .A(w_10_), .B(_395_), .C(_397_), .Y(_398_) );
INVX1 INVX1_569 ( .gnd(gnd), .vdd(vdd), .A(w_10_), .Y(_399_) );
INVX1 INVX1_570 ( .gnd(gnd), .vdd(vdd), .A(_395_), .Y(_400_) );
OAI21X1 OAI21X1_719 ( .gnd(gnd), .vdd(vdd), .A(_396_), .B(_400_), .C(_399_), .Y(_401_) );
AOI21X1 AOI21X1_91 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_401_), .C(_394_), .Y(_402_) );
NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_401_), .B(_398_), .Y(_403_) );
NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_403_), .Y(_404_) );
OAI22X1 OAI22X1_54 ( .gnd(gnd), .vdd(vdd), .A(_402_), .B(_404_), .C(_392_), .D(_386_), .Y(_405_) );
NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_385_), .Y(_406_) );
OAI21X1 OAI21X1_720 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf2), .B(_40__bF_buf1), .C(_406_), .Y(_407_) );
NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf2), .B(_391_), .Y(_408_) );
AOI21X1 AOI21X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf1), .B(_387_), .C(_408_), .Y(_409_) );
NAND3X1 NAND3X1_170 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_401_), .C(_398_), .Y(_410_) );
NOR3X1 NOR3X1_69 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_396_), .C(_400_), .Y(_411_) );
AOI21X1 AOI21X1_93 ( .gnd(gnd), .vdd(vdd), .A(_397_), .B(_395_), .C(w_10_), .Y(_412_) );
OAI21X1 OAI21X1_721 ( .gnd(gnd), .vdd(vdd), .A(_411_), .B(_412_), .C(_394_), .Y(_413_) );
NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_413_), .Y(_414_) );
NAND3X1 NAND3X1_171 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_407_), .C(_414_), .Y(_415_) );
NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_415_), .Y(_416_) );
OAI21X1 OAI21X1_722 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_350_), .C(_416_), .Y(_417_) );
AOI21X1 AOI21X1_94 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_336_), .C(_378_), .Y(_418_) );
NAND3X1 NAND3X1_172 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_415_), .C(_418_), .Y(_419_) );
AOI21X1 AOI21X1_95 ( .gnd(gnd), .vdd(vdd), .A(_417_), .B(_419_), .C(_3405__bF_buf4), .Y(_420_) );
OAI21X1 OAI21X1_723 ( .gnd(gnd), .vdd(vdd), .A(_343_), .B(_342_), .C(_332_), .Y(_421_) );
NAND3X1 NAND3X1_173 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_415_), .C(_421_), .Y(_422_) );
NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_416_), .Y(_423_) );
AOI21X1 AOI21X1_96 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_422_), .C(_3451__bF_buf0), .Y(_424_) );
OAI21X1 OAI21X1_724 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_420_), .C(_377_), .Y(_425_) );
NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_344_), .Y(_426_) );
NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_426_), .Y(_427_) );
AOI21X1 AOI21X1_97 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf0), .B(_352_), .C(_427_), .Y(_428_) );
NAND3X1 NAND3X1_174 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf4), .B(_422_), .C(_423_), .Y(_429_) );
NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_418_), .B(_416_), .Y(_430_) );
AOI21X1 AOI21X1_98 ( .gnd(gnd), .vdd(vdd), .A(_405_), .B(_415_), .C(_421_), .Y(_431_) );
OAI21X1 OAI21X1_725 ( .gnd(gnd), .vdd(vdd), .A(_431_), .B(_430_), .C(_3405__bF_buf3), .Y(_432_) );
NAND3X1 NAND3X1_175 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_432_), .C(_428_), .Y(_433_) );
NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(_425_), .B(_433_), .Y(_434_) );
AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_434_), .Y(_435_) );
NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_435_), .Y(_436_) );
OAI21X1 OAI21X1_726 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_434_), .C(_436_), .Y(_437_) );
INVX1 INVX1_571 ( .gnd(gnd), .vdd(vdd), .A(_3667__138_), .Y(_438_) );
NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_3432__bF_buf2), .Y(_439_) );
AOI22X1 AOI22X1_631 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_3433__bF_buf1), .C(a_reg_10_), .D(_113__bF_buf1), .Y(_440_) );
NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_440_), .B(_437_), .Y(_5__10_) );
NAND3X1 NAND3X1_176 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(_377_), .C(_432_), .Y(_441_) );
INVX1 INVX1_572 ( .gnd(gnd), .vdd(vdd), .A(_441_), .Y(_442_) );
NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(_442_), .B(_435_), .Y(_443_) );
OAI21X1 OAI21X1_727 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf2), .B(_431_), .C(_422_), .Y(_444_) );
AOI21X1 AOI21X1_99 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf1), .B(_406_), .C(_392_), .Y(_445_) );
OAI21X1 OAI21X1_728 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_445_), .C(_410_), .Y(_446_) );
NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(c_reg_11_), .B(b_reg_11_), .Y(_447_) );
INVX1 INVX1_573 ( .gnd(gnd), .vdd(vdd), .A(_447_), .Y(_448_) );
NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(c_reg_11_), .B(b_reg_11_), .Y(_449_) );
OAI21X1 OAI21X1_729 ( .gnd(gnd), .vdd(vdd), .A(_449_), .B(_448_), .C(d_reg_11_), .Y(_450_) );
INVX2 INVX2_26 ( .gnd(gnd), .vdd(vdd), .A(d_reg_11_), .Y(_451_) );
INVX1 INVX1_574 ( .gnd(gnd), .vdd(vdd), .A(_449_), .Y(_452_) );
NAND3X1 NAND3X1_177 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_447_), .C(_452_), .Y(_453_) );
NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_450_), .B(_453_), .Y(_454_) );
OAI21X1 OAI21X1_730 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf1), .B(_40__bF_buf3), .C(_454_), .Y(_455_) );
AOI21X1 AOI21X1_100 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_447_), .C(_449_), .Y(_456_) );
INVX1 INVX1_575 ( .gnd(gnd), .vdd(vdd), .A(c_reg_11_), .Y(_457_) );
NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(b_reg_11_), .B(_457_), .Y(_458_) );
OAI21X1 OAI21X1_731 ( .gnd(gnd), .vdd(vdd), .A(b_reg_11_), .B(d_reg_11_), .C(_458_), .Y(_459_) );
NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf1), .B(_459_), .Y(_460_) );
AOI21X1 AOI21X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf3), .B(_456_), .C(_460_), .Y(_461_) );
OAI21X1 OAI21X1_732 ( .gnd(gnd), .vdd(vdd), .A(_399_), .B(_396_), .C(_395_), .Y(_462_) );
NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(a_reg_6_), .B(e_reg_11_), .Y(_463_) );
NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(a_reg_6_), .B(e_reg_11_), .Y(_464_) );
INVX1 INVX1_576 ( .gnd(gnd), .vdd(vdd), .A(_464_), .Y(_465_) );
NAND3X1 NAND3X1_178 ( .gnd(gnd), .vdd(vdd), .A(w_11_), .B(_463_), .C(_465_), .Y(_466_) );
INVX1 INVX1_577 ( .gnd(gnd), .vdd(vdd), .A(w_11_), .Y(_467_) );
INVX1 INVX1_578 ( .gnd(gnd), .vdd(vdd), .A(_463_), .Y(_468_) );
OAI21X1 OAI21X1_733 ( .gnd(gnd), .vdd(vdd), .A(_464_), .B(_468_), .C(_467_), .Y(_469_) );
NAND3X1 NAND3X1_179 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_469_), .C(_466_), .Y(_470_) );
INVX1 INVX1_579 ( .gnd(gnd), .vdd(vdd), .A(_462_), .Y(_471_) );
NOR3X1 NOR3X1_70 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_464_), .C(_468_), .Y(_472_) );
AOI21X1 AOI21X1_102 ( .gnd(gnd), .vdd(vdd), .A(_465_), .B(_463_), .C(w_11_), .Y(_473_) );
OAI21X1 OAI21X1_734 ( .gnd(gnd), .vdd(vdd), .A(_472_), .B(_473_), .C(_471_), .Y(_474_) );
NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_470_), .B(_474_), .Y(_475_) );
AOI21X1 AOI21X1_103 ( .gnd(gnd), .vdd(vdd), .A(_455_), .B(_461_), .C(_475_), .Y(_476_) );
AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_453_), .B(_450_), .Y(_477_) );
OAI21X1 OAI21X1_735 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf4), .B(_477_), .C(_461_), .Y(_478_) );
AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_474_), .B(_470_), .Y(_479_) );
NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_478_), .Y(_480_) );
OAI21X1 OAI21X1_736 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_480_), .C(_446_), .Y(_481_) );
AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_385_), .B(_382_), .Y(_482_) );
OAI21X1 OAI21X1_737 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf3), .B(_482_), .C(_409_), .Y(_483_) );
INVX1 INVX1_580 ( .gnd(gnd), .vdd(vdd), .A(_410_), .Y(_484_) );
AOI21X1 AOI21X1_104 ( .gnd(gnd), .vdd(vdd), .A(_483_), .B(_413_), .C(_484_), .Y(_485_) );
NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(_479_), .B(_478_), .Y(_486_) );
NAND3X1 NAND3X1_180 ( .gnd(gnd), .vdd(vdd), .A(_461_), .B(_455_), .C(_475_), .Y(_487_) );
NAND3X1 NAND3X1_181 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(_485_), .Y(_488_) );
AOI22X1 AOI22X1_632 ( .gnd(gnd), .vdd(vdd), .A(_3448_), .B(_3450_), .C(_488_), .D(_481_), .Y(_489_) );
OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_3378_), .B(_3389_), .Y(_490_) );
NAND3X1 NAND3X1_182 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(_446_), .Y(_491_) );
OAI21X1 OAI21X1_738 ( .gnd(gnd), .vdd(vdd), .A(_476_), .B(_480_), .C(_485_), .Y(_492_) );
AOI22X1 AOI22X1_633 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_490_), .C(_492_), .D(_491_), .Y(_493_) );
OAI21X1 OAI21X1_739 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_493_), .C(_444_), .Y(_494_) );
AOI21X1 AOI21X1_105 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf2), .B(_423_), .C(_430_), .Y(_495_) );
NAND3X1 NAND3X1_183 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_492_), .C(_491_), .Y(_496_) );
NAND3X1 NAND3X1_184 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf0), .B(_488_), .C(_481_), .Y(_497_) );
NAND3X1 NAND3X1_185 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_496_), .C(_495_), .Y(_498_) );
NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_498_), .B(_494_), .Y(_499_) );
INVX1 INVX1_581 ( .gnd(gnd), .vdd(vdd), .A(_499_), .Y(_500_) );
AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_500_), .Y(_501_) );
OAI21X1 OAI21X1_740 ( .gnd(gnd), .vdd(vdd), .A(_500_), .B(_443_), .C(round_ctr_inc_bF_buf0), .Y(_502_) );
INVX1 INVX1_582 ( .gnd(gnd), .vdd(vdd), .A(_3667__139_), .Y(_503_) );
NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_3432__bF_buf1), .Y(_504_) );
AOI22X1 AOI22X1_634 ( .gnd(gnd), .vdd(vdd), .A(_504_), .B(_3433__bF_buf0), .C(a_reg_11_), .D(_113__bF_buf0), .Y(_505_) );
OAI21X1 OAI21X1_741 ( .gnd(gnd), .vdd(vdd), .A(_501_), .B(_502_), .C(_505_), .Y(_5__11_) );
AOI22X1 AOI22X1_635 ( .gnd(gnd), .vdd(vdd), .A(_494_), .B(_498_), .C(_425_), .D(_433_), .Y(_506_) );
NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_506_), .B(_369_), .Y(_507_) );
OAI21X1 OAI21X1_742 ( .gnd(gnd), .vdd(vdd), .A(_489_), .B(_493_), .C(_495_), .Y(_508_) );
NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_497_), .B(_496_), .Y(_509_) );
OAI21X1 OAI21X1_743 ( .gnd(gnd), .vdd(vdd), .A(_495_), .B(_509_), .C(_441_), .Y(_510_) );
AOI22X1 AOI22X1_636 ( .gnd(gnd), .vdd(vdd), .A(_508_), .B(_510_), .C(_373_), .D(_506_), .Y(_511_) );
OAI21X1 OAI21X1_744 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_242_), .C(_511_), .Y(_512_) );
AOI21X1 AOI21X1_106 ( .gnd(gnd), .vdd(vdd), .A(_486_), .B(_487_), .C(_446_), .Y(_513_) );
OAI21X1 OAI21X1_745 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf3), .B(_513_), .C(_491_), .Y(_514_) );
NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(_456_), .B(_3451__bF_buf1), .Y(_515_) );
OAI21X1 OAI21X1_746 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf0), .B(_459_), .C(_515_), .Y(_516_) );
AOI21X1 AOI21X1_107 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf0), .B(_454_), .C(_516_), .Y(_517_) );
OAI21X1 OAI21X1_747 ( .gnd(gnd), .vdd(vdd), .A(_475_), .B(_517_), .C(_470_), .Y(_518_) );
INVX2 INVX2_27 ( .gnd(gnd), .vdd(vdd), .A(d_reg_12_), .Y(_519_) );
NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(c_reg_12_), .B(b_reg_12_), .Y(_520_) );
NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_520_), .Y(_521_) );
NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(c_reg_12_), .B(b_reg_12_), .Y(_522_) );
AOI21X1 AOI21X1_108 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_522_), .C(_520_), .Y(_523_) );
OAI21X1 OAI21X1_748 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_522_), .C(_523_), .Y(_524_) );
NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(_521_), .B(_524_), .Y(_525_) );
INVX1 INVX1_583 ( .gnd(gnd), .vdd(vdd), .A(c_reg_12_), .Y(_526_) );
NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(b_reg_12_), .B(_526_), .Y(_527_) );
OAI21X1 OAI21X1_749 ( .gnd(gnd), .vdd(vdd), .A(b_reg_12_), .B(d_reg_12_), .C(_527_), .Y(_528_) );
NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf4), .B(_528_), .Y(_529_) );
AOI21X1 AOI21X1_109 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf0), .B(_523_), .C(_529_), .Y(_530_) );
OAI21X1 OAI21X1_750 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf2), .B(_525_), .C(_530_), .Y(_531_) );
OAI21X1 OAI21X1_751 ( .gnd(gnd), .vdd(vdd), .A(_467_), .B(_464_), .C(_463_), .Y(_532_) );
NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(a_reg_7_), .B(e_reg_12_), .Y(_533_) );
NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(a_reg_7_), .B(e_reg_12_), .Y(_534_) );
INVX1 INVX1_584 ( .gnd(gnd), .vdd(vdd), .A(_534_), .Y(_535_) );
NAND3X1 NAND3X1_186 ( .gnd(gnd), .vdd(vdd), .A(w_12_), .B(_533_), .C(_535_), .Y(_536_) );
INVX1 INVX1_585 ( .gnd(gnd), .vdd(vdd), .A(w_12_), .Y(_537_) );
INVX1 INVX1_586 ( .gnd(gnd), .vdd(vdd), .A(_533_), .Y(_538_) );
OAI21X1 OAI21X1_752 ( .gnd(gnd), .vdd(vdd), .A(_534_), .B(_538_), .C(_537_), .Y(_539_) );
NAND3X1 NAND3X1_187 ( .gnd(gnd), .vdd(vdd), .A(_532_), .B(_539_), .C(_536_), .Y(_540_) );
NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_539_), .B(_536_), .Y(_541_) );
NAND3X1 NAND3X1_188 ( .gnd(gnd), .vdd(vdd), .A(_463_), .B(_466_), .C(_541_), .Y(_542_) );
NAND3X1 NAND3X1_189 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_542_), .C(_531_), .Y(_543_) );
INVX1 INVX1_587 ( .gnd(gnd), .vdd(vdd), .A(_525_), .Y(_544_) );
NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(_523_), .B(_3451__bF_buf4), .Y(_545_) );
OAI21X1 OAI21X1_753 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf3), .B(_528_), .C(_545_), .Y(_546_) );
AOI21X1 AOI21X1_110 ( .gnd(gnd), .vdd(vdd), .A(_544_), .B(_3474__bF_buf4), .C(_546_), .Y(_547_) );
NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_542_), .Y(_548_) );
NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_547_), .Y(_549_) );
NAND3X1 NAND3X1_190 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_549_), .C(_518_), .Y(_550_) );
INVX1 INVX1_588 ( .gnd(gnd), .vdd(vdd), .A(_470_), .Y(_551_) );
AOI21X1 AOI21X1_111 ( .gnd(gnd), .vdd(vdd), .A(_478_), .B(_474_), .C(_551_), .Y(_552_) );
OAI21X1 OAI21X1_754 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf2), .B(_40__bF_buf2), .C(_544_), .Y(_553_) );
AOI21X1 AOI21X1_112 ( .gnd(gnd), .vdd(vdd), .A(_553_), .B(_530_), .C(_548_), .Y(_554_) );
AOI21X1 AOI21X1_113 ( .gnd(gnd), .vdd(vdd), .A(_540_), .B(_542_), .C(_531_), .Y(_555_) );
OAI21X1 OAI21X1_755 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_554_), .C(_552_), .Y(_556_) );
AOI21X1 AOI21X1_114 ( .gnd(gnd), .vdd(vdd), .A(_556_), .B(_550_), .C(_3406__bF_buf1), .Y(_557_) );
OAI21X1 OAI21X1_756 ( .gnd(gnd), .vdd(vdd), .A(_555_), .B(_554_), .C(_518_), .Y(_558_) );
NAND3X1 NAND3X1_191 ( .gnd(gnd), .vdd(vdd), .A(_543_), .B(_552_), .C(_549_), .Y(_559_) );
AOI21X1 AOI21X1_115 ( .gnd(gnd), .vdd(vdd), .A(_558_), .B(_559_), .C(_3474__bF_buf3), .Y(_560_) );
OAI21X1 OAI21X1_757 ( .gnd(gnd), .vdd(vdd), .A(_560_), .B(_557_), .C(_514_), .Y(_561_) );
NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_487_), .B(_486_), .Y(_562_) );
NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_485_), .B(_562_), .Y(_563_) );
AOI21X1 AOI21X1_116 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_492_), .C(_563_), .Y(_564_) );
NAND3X1 NAND3X1_192 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf2), .B(_559_), .C(_558_), .Y(_565_) );
NAND3X1 NAND3X1_193 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf0), .B(_550_), .C(_556_), .Y(_566_) );
NAND3X1 NAND3X1_194 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_566_), .C(_564_), .Y(_567_) );
NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_567_), .B(_561_), .Y(_568_) );
XNOR2X1 XNOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_568_), .Y(_569_) );
INVX1 INVX1_589 ( .gnd(gnd), .vdd(vdd), .A(_3667__140_), .Y(_570_) );
NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_3432__bF_buf0), .Y(_571_) );
AOI22X1 AOI22X1_637 ( .gnd(gnd), .vdd(vdd), .A(_571_), .B(_3433__bF_buf11), .C(a_reg_12_), .D(_113__bF_buf4), .Y(_572_) );
OAI21X1 OAI21X1_758 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_569_), .C(_572_), .Y(_5__12_) );
AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_512_), .B(_568_), .Y(_573_) );
NAND3X1 NAND3X1_195 ( .gnd(gnd), .vdd(vdd), .A(_565_), .B(_566_), .C(_514_), .Y(_574_) );
AOI21X1 AOI21X1_117 ( .gnd(gnd), .vdd(vdd), .A(_549_), .B(_543_), .C(_518_), .Y(_575_) );
OAI21X1 OAI21X1_759 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf1), .B(_575_), .C(_550_), .Y(_576_) );
INVX1 INVX1_590 ( .gnd(gnd), .vdd(vdd), .A(_540_), .Y(_577_) );
NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(c_reg_13_), .B(b_reg_13_), .Y(_578_) );
INVX1 INVX1_591 ( .gnd(gnd), .vdd(vdd), .A(_578_), .Y(_579_) );
NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(c_reg_13_), .B(b_reg_13_), .Y(_580_) );
OAI21X1 OAI21X1_760 ( .gnd(gnd), .vdd(vdd), .A(_580_), .B(_579_), .C(d_reg_13_), .Y(_581_) );
INVX2 INVX2_28 ( .gnd(gnd), .vdd(vdd), .A(d_reg_13_), .Y(_582_) );
INVX1 INVX1_592 ( .gnd(gnd), .vdd(vdd), .A(_580_), .Y(_583_) );
NAND3X1 NAND3X1_196 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_578_), .C(_583_), .Y(_584_) );
NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_581_), .B(_584_), .Y(_585_) );
INVX1 INVX1_593 ( .gnd(gnd), .vdd(vdd), .A(_585_), .Y(_586_) );
AOI21X1 AOI21X1_118 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_578_), .C(_580_), .Y(_587_) );
INVX1 INVX1_594 ( .gnd(gnd), .vdd(vdd), .A(c_reg_13_), .Y(_588_) );
NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(b_reg_13_), .B(_588_), .Y(_589_) );
OAI21X1 OAI21X1_761 ( .gnd(gnd), .vdd(vdd), .A(b_reg_13_), .B(d_reg_13_), .C(_589_), .Y(_590_) );
NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf2), .B(_590_), .Y(_591_) );
AOI21X1 AOI21X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf3), .B(_587_), .C(_591_), .Y(_592_) );
OAI21X1 OAI21X1_762 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf4), .B(_586_), .C(_592_), .Y(_593_) );
OAI21X1 OAI21X1_763 ( .gnd(gnd), .vdd(vdd), .A(_537_), .B(_534_), .C(_533_), .Y(_594_) );
INVX1 INVX1_595 ( .gnd(gnd), .vdd(vdd), .A(_594_), .Y(_595_) );
NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(a_reg_8_), .B(e_reg_13_), .Y(_596_) );
NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(a_reg_8_), .B(e_reg_13_), .Y(_597_) );
INVX1 INVX1_596 ( .gnd(gnd), .vdd(vdd), .A(_597_), .Y(_598_) );
NAND3X1 NAND3X1_197 ( .gnd(gnd), .vdd(vdd), .A(w_13_), .B(_596_), .C(_598_), .Y(_599_) );
INVX1 INVX1_597 ( .gnd(gnd), .vdd(vdd), .A(w_13_), .Y(_600_) );
INVX1 INVX1_598 ( .gnd(gnd), .vdd(vdd), .A(_596_), .Y(_601_) );
OAI21X1 OAI21X1_764 ( .gnd(gnd), .vdd(vdd), .A(_597_), .B(_601_), .C(_600_), .Y(_602_) );
AOI21X1 AOI21X1_120 ( .gnd(gnd), .vdd(vdd), .A(_599_), .B(_602_), .C(_595_), .Y(_603_) );
NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_602_), .B(_599_), .Y(_604_) );
NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_604_), .Y(_605_) );
OAI21X1 OAI21X1_765 ( .gnd(gnd), .vdd(vdd), .A(_603_), .B(_605_), .C(_593_), .Y(_606_) );
OAI21X1 OAI21X1_766 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf1), .B(_40__bF_buf1), .C(_585_), .Y(_607_) );
NAND3X1 NAND3X1_198 ( .gnd(gnd), .vdd(vdd), .A(_594_), .B(_602_), .C(_599_), .Y(_608_) );
NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_595_), .B(_604_), .Y(_609_) );
NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(_608_), .B(_609_), .Y(_610_) );
NAND3X1 NAND3X1_199 ( .gnd(gnd), .vdd(vdd), .A(_607_), .B(_592_), .C(_610_), .Y(_611_) );
NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_611_), .B(_606_), .Y(_612_) );
OAI21X1 OAI21X1_767 ( .gnd(gnd), .vdd(vdd), .A(_577_), .B(_554_), .C(_612_), .Y(_613_) );
AOI21X1 AOI21X1_121 ( .gnd(gnd), .vdd(vdd), .A(_531_), .B(_542_), .C(_577_), .Y(_614_) );
NAND3X1 NAND3X1_200 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_611_), .C(_614_), .Y(_615_) );
NAND3X1 NAND3X1_201 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf0), .B(_615_), .C(_613_), .Y(_616_) );
OAI21X1 OAI21X1_768 ( .gnd(gnd), .vdd(vdd), .A(_548_), .B(_547_), .C(_540_), .Y(_617_) );
NAND3X1 NAND3X1_202 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_611_), .C(_617_), .Y(_618_) );
NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_612_), .Y(_619_) );
NAND3X1 NAND3X1_203 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_618_), .C(_619_), .Y(_620_) );
NAND3X1 NAND3X1_204 ( .gnd(gnd), .vdd(vdd), .A(_576_), .B(_620_), .C(_616_), .Y(_621_) );
INVX1 INVX1_599 ( .gnd(gnd), .vdd(vdd), .A(_621_), .Y(_622_) );
AOI21X1 AOI21X1_122 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_620_), .C(_576_), .Y(_623_) );
OAI21X1 OAI21X1_769 ( .gnd(gnd), .vdd(vdd), .A(_623_), .B(_622_), .C(_574_), .Y(_624_) );
INVX1 INVX1_600 ( .gnd(gnd), .vdd(vdd), .A(_574_), .Y(_625_) );
AOI21X1 AOI21X1_123 ( .gnd(gnd), .vdd(vdd), .A(_619_), .B(_618_), .C(_3472_), .Y(_626_) );
AOI22X1 AOI22X1_638 ( .gnd(gnd), .vdd(vdd), .A(_3448_), .B(_3450_), .C(_615_), .D(_613_), .Y(_627_) );
OAI21X1 OAI21X1_770 ( .gnd(gnd), .vdd(vdd), .A(_627_), .B(_626_), .C(_576_), .Y(_628_) );
INVX1 INVX1_601 ( .gnd(gnd), .vdd(vdd), .A(_550_), .Y(_629_) );
AOI21X1 AOI21X1_124 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf3), .B(_556_), .C(_629_), .Y(_630_) );
NAND3X1 NAND3X1_205 ( .gnd(gnd), .vdd(vdd), .A(_616_), .B(_620_), .C(_630_), .Y(_631_) );
NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_631_), .B(_628_), .Y(_632_) );
OAI21X1 OAI21X1_771 ( .gnd(gnd), .vdd(vdd), .A(_625_), .B(_573_), .C(_632_), .Y(_633_) );
OAI21X1 OAI21X1_772 ( .gnd(gnd), .vdd(vdd), .A(_573_), .B(_624_), .C(_633_), .Y(_634_) );
INVX1 INVX1_602 ( .gnd(gnd), .vdd(vdd), .A(_3667__141_), .Y(_635_) );
OAI21X1 OAI21X1_773 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_635_), .Y(_636_) );
AOI22X1 AOI22X1_639 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf10), .B(_636_), .C(a_reg_13_), .D(_113__bF_buf3), .Y(_637_) );
OAI21X1 OAI21X1_774 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_634_), .C(_637_), .Y(_5__13_) );
AOI22X1 AOI22X1_640 ( .gnd(gnd), .vdd(vdd), .A(_561_), .B(_567_), .C(_631_), .D(_628_), .Y(_638_) );
NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_512_), .Y(_639_) );
OAI21X1 OAI21X1_775 ( .gnd(gnd), .vdd(vdd), .A(_574_), .B(_623_), .C(_621_), .Y(_640_) );
INVX1 INVX1_603 ( .gnd(gnd), .vdd(vdd), .A(_640_), .Y(_641_) );
NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_641_), .B(_639_), .Y(_642_) );
AOI21X1 AOI21X1_125 ( .gnd(gnd), .vdd(vdd), .A(_606_), .B(_611_), .C(_617_), .Y(_643_) );
OAI21X1 OAI21X1_776 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf3), .B(_643_), .C(_618_), .Y(_644_) );
NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_587_), .B(_3451__bF_buf2), .Y(_645_) );
OAI21X1 OAI21X1_777 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf1), .B(_590_), .C(_645_), .Y(_646_) );
AOI21X1 AOI21X1_126 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf0), .B(_585_), .C(_646_), .Y(_647_) );
OAI21X1 OAI21X1_778 ( .gnd(gnd), .vdd(vdd), .A(_610_), .B(_647_), .C(_608_), .Y(_648_) );
NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(c_reg_14_), .B(b_reg_14_), .Y(_649_) );
NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(c_reg_14_), .B(b_reg_14_), .Y(_650_) );
INVX1 INVX1_604 ( .gnd(gnd), .vdd(vdd), .A(_650_), .Y(_651_) );
NAND3X1 NAND3X1_206 ( .gnd(gnd), .vdd(vdd), .A(d_reg_14_), .B(_649_), .C(_651_), .Y(_652_) );
INVX2 INVX2_29 ( .gnd(gnd), .vdd(vdd), .A(d_reg_14_), .Y(_653_) );
INVX1 INVX1_605 ( .gnd(gnd), .vdd(vdd), .A(_649_), .Y(_654_) );
OAI21X1 OAI21X1_779 ( .gnd(gnd), .vdd(vdd), .A(_650_), .B(_654_), .C(_653_), .Y(_655_) );
NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(_655_), .B(_652_), .Y(_656_) );
AOI21X1 AOI21X1_127 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_649_), .C(_650_), .Y(_657_) );
OAI21X1 OAI21X1_780 ( .gnd(gnd), .vdd(vdd), .A(b_reg_14_), .B(_653_), .C(_649_), .Y(_658_) );
AOI22X1 AOI22X1_641 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf3), .B(_658_), .C(_3451__bF_buf1), .D(_657_), .Y(_659_) );
OAI21X1 OAI21X1_781 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf2), .B(_656_), .C(_659_), .Y(_660_) );
OAI21X1 OAI21X1_782 ( .gnd(gnd), .vdd(vdd), .A(_600_), .B(_597_), .C(_596_), .Y(_661_) );
NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(a_reg_9_), .B(e_reg_14_), .Y(_662_) );
NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(a_reg_9_), .B(e_reg_14_), .Y(_663_) );
INVX1 INVX1_606 ( .gnd(gnd), .vdd(vdd), .A(_663_), .Y(_664_) );
NAND3X1 NAND3X1_207 ( .gnd(gnd), .vdd(vdd), .A(w_14_), .B(_662_), .C(_664_), .Y(_665_) );
INVX1 INVX1_607 ( .gnd(gnd), .vdd(vdd), .A(w_14_), .Y(_666_) );
INVX1 INVX1_608 ( .gnd(gnd), .vdd(vdd), .A(_662_), .Y(_667_) );
OAI21X1 OAI21X1_783 ( .gnd(gnd), .vdd(vdd), .A(_663_), .B(_667_), .C(_666_), .Y(_668_) );
NAND3X1 NAND3X1_208 ( .gnd(gnd), .vdd(vdd), .A(_661_), .B(_668_), .C(_665_), .Y(_669_) );
NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_668_), .B(_665_), .Y(_670_) );
NAND3X1 NAND3X1_209 ( .gnd(gnd), .vdd(vdd), .A(_596_), .B(_599_), .C(_670_), .Y(_671_) );
NAND3X1 NAND3X1_210 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_671_), .C(_660_), .Y(_672_) );
INVX1 INVX1_609 ( .gnd(gnd), .vdd(vdd), .A(_656_), .Y(_673_) );
INVX1 INVX1_610 ( .gnd(gnd), .vdd(vdd), .A(_657_), .Y(_674_) );
NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(_658_), .B(_3447__bF_buf2), .Y(_675_) );
OAI21X1 OAI21X1_784 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf1), .B(_674_), .C(_675_), .Y(_676_) );
AOI21X1 AOI21X1_128 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf4), .B(_673_), .C(_676_), .Y(_677_) );
NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_671_), .Y(_678_) );
NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_677_), .Y(_679_) );
NAND3X1 NAND3X1_211 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_679_), .C(_648_), .Y(_680_) );
INVX1 INVX1_611 ( .gnd(gnd), .vdd(vdd), .A(_608_), .Y(_681_) );
AOI21X1 AOI21X1_129 ( .gnd(gnd), .vdd(vdd), .A(_593_), .B(_609_), .C(_681_), .Y(_682_) );
INVX1 INVX1_612 ( .gnd(gnd), .vdd(vdd), .A(_672_), .Y(_683_) );
AOI21X1 AOI21X1_130 ( .gnd(gnd), .vdd(vdd), .A(_669_), .B(_671_), .C(_660_), .Y(_684_) );
OAI21X1 OAI21X1_785 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_683_), .C(_682_), .Y(_685_) );
AOI21X1 AOI21X1_131 ( .gnd(gnd), .vdd(vdd), .A(_685_), .B(_680_), .C(_3405__bF_buf0), .Y(_686_) );
OAI21X1 OAI21X1_786 ( .gnd(gnd), .vdd(vdd), .A(_684_), .B(_683_), .C(_648_), .Y(_687_) );
NAND3X1 NAND3X1_212 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_679_), .C(_682_), .Y(_688_) );
AOI21X1 AOI21X1_132 ( .gnd(gnd), .vdd(vdd), .A(_687_), .B(_688_), .C(_3451__bF_buf0), .Y(_689_) );
OAI21X1 OAI21X1_787 ( .gnd(gnd), .vdd(vdd), .A(_689_), .B(_686_), .C(_644_), .Y(_690_) );
NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_614_), .B(_612_), .Y(_691_) );
AOI21X1 AOI21X1_133 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_619_), .C(_691_), .Y(_692_) );
NAND3X1 NAND3X1_213 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf4), .B(_688_), .C(_687_), .Y(_693_) );
NAND3X1 NAND3X1_214 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf5), .B(_680_), .C(_685_), .Y(_694_) );
NAND3X1 NAND3X1_215 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_694_), .C(_692_), .Y(_695_) );
NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_695_), .B(_690_), .Y(_696_) );
AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_642_), .B(_696_), .Y(_697_) );
OAI21X1 OAI21X1_788 ( .gnd(gnd), .vdd(vdd), .A(_696_), .B(_642_), .C(round_ctr_inc_bF_buf11), .Y(_698_) );
INVX2 INVX2_30 ( .gnd(gnd), .vdd(vdd), .A(_3667__142_), .Y(_699_) );
NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_3432__bF_buf11), .Y(_700_) );
AOI22X1 AOI22X1_642 ( .gnd(gnd), .vdd(vdd), .A(_700_), .B(_3433__bF_buf9), .C(a_reg_14_), .D(_113__bF_buf2), .Y(_701_) );
OAI21X1 OAI21X1_789 ( .gnd(gnd), .vdd(vdd), .A(_697_), .B(_698_), .C(_701_), .Y(_5__14_) );
NAND3X1 NAND3X1_216 ( .gnd(gnd), .vdd(vdd), .A(_693_), .B(_694_), .C(_644_), .Y(_702_) );
INVX1 INVX1_613 ( .gnd(gnd), .vdd(vdd), .A(_702_), .Y(_703_) );
NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(_703_), .B(_697_), .Y(_704_) );
AOI21X1 AOI21X1_134 ( .gnd(gnd), .vdd(vdd), .A(_672_), .B(_679_), .C(_648_), .Y(_705_) );
OAI21X1 OAI21X1_790 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf3), .B(_705_), .C(_680_), .Y(_706_) );
INVX1 INVX1_614 ( .gnd(gnd), .vdd(vdd), .A(_669_), .Y(_707_) );
AOI21X1 AOI21X1_135 ( .gnd(gnd), .vdd(vdd), .A(_660_), .B(_671_), .C(_707_), .Y(_708_) );
INVX2 INVX2_31 ( .gnd(gnd), .vdd(vdd), .A(b_reg_15_), .Y(_709_) );
AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(c_reg_15_), .B(b_reg_15_), .Y(_710_) );
AOI21X1 AOI21X1_136 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(d_reg_15_), .C(_710_), .Y(_711_) );
NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_711_), .B(_3447__bF_buf1), .Y(_712_) );
NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(c_reg_15_), .B(b_reg_15_), .Y(_713_) );
OAI21X1 OAI21X1_791 ( .gnd(gnd), .vdd(vdd), .A(c_reg_15_), .B(b_reg_15_), .C(d_reg_15_), .Y(_714_) );
NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_713_), .B(_714_), .Y(_715_) );
NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(_715_), .B(_3451__bF_buf2), .Y(_716_) );
INVX1 INVX1_615 ( .gnd(gnd), .vdd(vdd), .A(_3402_), .Y(_717_) );
INVX2 INVX2_32 ( .gnd(gnd), .vdd(vdd), .A(d_reg_15_), .Y(_718_) );
NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(c_reg_15_), .B(b_reg_15_), .Y(_719_) );
NAND3X1 NAND3X1_217 ( .gnd(gnd), .vdd(vdd), .A(c_reg_15_), .B(b_reg_15_), .C(d_reg_15_), .Y(_720_) );
AOI22X1 AOI22X1_643 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_719_), .C(_720_), .D(_715_), .Y(_721_) );
AOI22X1 AOI22X1_644 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_717_), .C(_3405__bF_buf4), .D(_721_), .Y(_722_) );
NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_716_), .B(_722_), .Y(_723_) );
OAI21X1 OAI21X1_792 ( .gnd(gnd), .vdd(vdd), .A(_666_), .B(_663_), .C(_662_), .Y(_724_) );
NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(a_reg_10_), .B(e_reg_15_), .Y(_725_) );
NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(a_reg_10_), .B(e_reg_15_), .Y(_726_) );
INVX1 INVX1_616 ( .gnd(gnd), .vdd(vdd), .A(_726_), .Y(_727_) );
NAND3X1 NAND3X1_218 ( .gnd(gnd), .vdd(vdd), .A(w_15_), .B(_725_), .C(_727_), .Y(_728_) );
INVX1 INVX1_617 ( .gnd(gnd), .vdd(vdd), .A(w_15_), .Y(_729_) );
AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(a_reg_10_), .B(e_reg_15_), .Y(_730_) );
OAI21X1 OAI21X1_793 ( .gnd(gnd), .vdd(vdd), .A(_726_), .B(_730_), .C(_729_), .Y(_731_) );
NAND3X1 NAND3X1_219 ( .gnd(gnd), .vdd(vdd), .A(_724_), .B(_731_), .C(_728_), .Y(_732_) );
INVX1 INVX1_618 ( .gnd(gnd), .vdd(vdd), .A(_724_), .Y(_733_) );
NOR3X1 NOR3X1_71 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_726_), .C(_730_), .Y(_734_) );
AOI21X1 AOI21X1_137 ( .gnd(gnd), .vdd(vdd), .A(_727_), .B(_725_), .C(w_15_), .Y(_735_) );
OAI21X1 OAI21X1_794 ( .gnd(gnd), .vdd(vdd), .A(_734_), .B(_735_), .C(_733_), .Y(_736_) );
AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_736_), .B(_732_), .Y(_737_) );
AOI21X1 AOI21X1_138 ( .gnd(gnd), .vdd(vdd), .A(_723_), .B(_712_), .C(_737_), .Y(_738_) );
AOI22X1 AOI22X1_645 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf0), .B(_711_), .C(_716_), .D(_722_), .Y(_739_) );
AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_739_), .B(_737_), .Y(_740_) );
OAI21X1 OAI21X1_795 ( .gnd(gnd), .vdd(vdd), .A(_738_), .B(_740_), .C(_708_), .Y(_741_) );
OAI21X1 OAI21X1_796 ( .gnd(gnd), .vdd(vdd), .A(_678_), .B(_677_), .C(_669_), .Y(_742_) );
INVX1 INVX1_619 ( .gnd(gnd), .vdd(vdd), .A(_716_), .Y(_743_) );
INVX1 INVX1_620 ( .gnd(gnd), .vdd(vdd), .A(c_reg_15_), .Y(_744_) );
NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_709_), .Y(_745_) );
NAND3X1 NAND3X1_220 ( .gnd(gnd), .vdd(vdd), .A(d_reg_15_), .B(_713_), .C(_745_), .Y(_746_) );
OAI21X1 OAI21X1_797 ( .gnd(gnd), .vdd(vdd), .A(_719_), .B(_710_), .C(_718_), .Y(_747_) );
NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(_747_), .B(_746_), .Y(_748_) );
OAI21X1 OAI21X1_798 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf1), .B(_748_), .C(_3411__bF_buf0), .Y(_749_) );
OAI21X1 OAI21X1_799 ( .gnd(gnd), .vdd(vdd), .A(_743_), .B(_749_), .C(_712_), .Y(_750_) );
NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_736_), .Y(_751_) );
NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_750_), .Y(_752_) );
NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_737_), .B(_739_), .Y(_753_) );
NAND3X1 NAND3X1_221 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_753_), .C(_742_), .Y(_754_) );
AOI21X1 AOI21X1_139 ( .gnd(gnd), .vdd(vdd), .A(_741_), .B(_754_), .C(_3411__bF_buf4), .Y(_755_) );
AOI21X1 AOI21X1_140 ( .gnd(gnd), .vdd(vdd), .A(_752_), .B(_753_), .C(_742_), .Y(_756_) );
NOR3X1 NOR3X1_72 ( .gnd(gnd), .vdd(vdd), .A(_708_), .B(_738_), .C(_740_), .Y(_757_) );
NOR3X1 NOR3X1_73 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf4), .B(_756_), .C(_757_), .Y(_758_) );
OAI21X1 OAI21X1_800 ( .gnd(gnd), .vdd(vdd), .A(_755_), .B(_758_), .C(_706_), .Y(_759_) );
INVX1 INVX1_621 ( .gnd(gnd), .vdd(vdd), .A(_680_), .Y(_760_) );
AOI21X1 AOI21X1_141 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf3), .B(_685_), .C(_760_), .Y(_761_) );
OAI21X1 OAI21X1_801 ( .gnd(gnd), .vdd(vdd), .A(_756_), .B(_757_), .C(_3447__bF_buf3), .Y(_762_) );
NAND3X1 NAND3X1_222 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf3), .B(_754_), .C(_741_), .Y(_763_) );
NAND3X1 NAND3X1_223 ( .gnd(gnd), .vdd(vdd), .A(_763_), .B(_762_), .C(_761_), .Y(_764_) );
NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_764_), .B(_759_), .Y(_765_) );
INVX1 INVX1_622 ( .gnd(gnd), .vdd(vdd), .A(_765_), .Y(_766_) );
AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_704_), .B(_766_), .Y(_767_) );
OAI21X1 OAI21X1_802 ( .gnd(gnd), .vdd(vdd), .A(_766_), .B(_704_), .C(round_ctr_inc_bF_buf10), .Y(_768_) );
INVX1 INVX1_623 ( .gnd(gnd), .vdd(vdd), .A(_3667__143_), .Y(_769_) );
NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_3432__bF_buf10), .Y(_770_) );
AOI22X1 AOI22X1_646 ( .gnd(gnd), .vdd(vdd), .A(_770_), .B(_3433__bF_buf8), .C(a_reg_15_), .D(_113__bF_buf1), .Y(_771_) );
OAI21X1 OAI21X1_803 ( .gnd(gnd), .vdd(vdd), .A(_767_), .B(_768_), .C(_771_), .Y(_5__15_) );
NAND3X1 NAND3X1_224 ( .gnd(gnd), .vdd(vdd), .A(_121_), .B(_237_), .C(_120_), .Y(_772_) );
AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_369_), .B(_506_), .Y(_773_) );
AOI22X1 AOI22X1_647 ( .gnd(gnd), .vdd(vdd), .A(_690_), .B(_695_), .C(_764_), .D(_759_), .Y(_774_) );
NAND3X1 NAND3X1_225 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_774_), .C(_773_), .Y(_775_) );
AOI21X1 AOI21X1_142 ( .gnd(gnd), .vdd(vdd), .A(_772_), .B(_240_), .C(_775_), .Y(_776_) );
NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(_638_), .B(_774_), .Y(_777_) );
NAND3X1 NAND3X1_226 ( .gnd(gnd), .vdd(vdd), .A(_706_), .B(_763_), .C(_762_), .Y(_778_) );
AOI21X1 AOI21X1_143 ( .gnd(gnd), .vdd(vdd), .A(_762_), .B(_763_), .C(_706_), .Y(_779_) );
OAI21X1 OAI21X1_804 ( .gnd(gnd), .vdd(vdd), .A(_702_), .B(_779_), .C(_778_), .Y(_780_) );
AOI21X1 AOI21X1_144 ( .gnd(gnd), .vdd(vdd), .A(_774_), .B(_640_), .C(_780_), .Y(_781_) );
OAI21X1 OAI21X1_805 ( .gnd(gnd), .vdd(vdd), .A(_511_), .B(_777_), .C(_781_), .Y(_782_) );
OAI21X1 OAI21X1_806 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf2), .B(_756_), .C(_754_), .Y(_783_) );
INVX1 INVX1_624 ( .gnd(gnd), .vdd(vdd), .A(_783_), .Y(_784_) );
OAI21X1 OAI21X1_807 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3437__bF_buf2), .C(_3473_), .Y(_785_) );
INVX4 INVX4_5 ( .gnd(gnd), .vdd(vdd), .A(_785_), .Y(_786_) );
OAI21X1 OAI21X1_808 ( .gnd(gnd), .vdd(vdd), .A(_751_), .B(_750_), .C(_732_), .Y(_787_) );
INVX2 INVX2_33 ( .gnd(gnd), .vdd(vdd), .A(d_reg_16_), .Y(_788_) );
XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(c_reg_16_), .B(b_reg_16_), .Y(_789_) );
NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_789_), .Y(_790_) );
AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_789_), .B(_788_), .Y(_791_) );
OAI21X1 OAI21X1_809 ( .gnd(gnd), .vdd(vdd), .A(_790_), .B(_791_), .C(_3474__bF_buf3), .Y(_792_) );
INVX1 INVX1_625 ( .gnd(gnd), .vdd(vdd), .A(c_reg_16_), .Y(_793_) );
INVX2 INVX2_34 ( .gnd(gnd), .vdd(vdd), .A(b_reg_16_), .Y(_794_) );
OAI21X1 OAI21X1_810 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_794_), .C(_788_), .Y(_795_) );
OAI21X1 OAI21X1_811 ( .gnd(gnd), .vdd(vdd), .A(c_reg_16_), .B(b_reg_16_), .C(_795_), .Y(_796_) );
NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_796_), .B(_3405__bF_buf2), .Y(_797_) );
OAI21X1 OAI21X1_812 ( .gnd(gnd), .vdd(vdd), .A(c_reg_16_), .B(_794_), .C(_795_), .Y(_798_) );
NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf2), .B(_798_), .Y(_799_) );
NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_799_), .B(_797_), .Y(_800_) );
AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(_800_), .B(_792_), .Y(_801_) );
OAI21X1 OAI21X1_813 ( .gnd(gnd), .vdd(vdd), .A(_729_), .B(_726_), .C(_725_), .Y(_802_) );
INVX1 INVX1_626 ( .gnd(gnd), .vdd(vdd), .A(_802_), .Y(_803_) );
INVX1 INVX1_627 ( .gnd(gnd), .vdd(vdd), .A(w_16_), .Y(_804_) );
NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(a_reg_11_), .B(e_reg_16_), .Y(_805_) );
INVX1 INVX1_628 ( .gnd(gnd), .vdd(vdd), .A(a_reg_11_), .Y(_806_) );
INVX1 INVX1_629 ( .gnd(gnd), .vdd(vdd), .A(e_reg_16_), .Y(_807_) );
NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_806_), .B(_807_), .Y(_808_) );
NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_805_), .B(_808_), .Y(_809_) );
NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_804_), .B(_809_), .Y(_810_) );
AOI21X1 AOI21X1_145 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(_805_), .C(w_16_), .Y(_811_) );
OAI21X1 OAI21X1_814 ( .gnd(gnd), .vdd(vdd), .A(_811_), .B(_810_), .C(_803_), .Y(_812_) );
OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_809_), .B(_804_), .Y(_813_) );
INVX1 INVX1_630 ( .gnd(gnd), .vdd(vdd), .A(_811_), .Y(_814_) );
NAND3X1 NAND3X1_227 ( .gnd(gnd), .vdd(vdd), .A(_802_), .B(_814_), .C(_813_), .Y(_815_) );
NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_815_), .Y(_816_) );
NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_801_), .Y(_817_) );
NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_792_), .B(_800_), .Y(_818_) );
NAND3X1 NAND3X1_228 ( .gnd(gnd), .vdd(vdd), .A(_812_), .B(_815_), .C(_818_), .Y(_819_) );
NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(_819_), .B(_817_), .Y(_820_) );
NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_820_), .Y(_821_) );
XNOR2X1 XNOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_816_), .Y(_822_) );
NAND3X1 NAND3X1_229 ( .gnd(gnd), .vdd(vdd), .A(_732_), .B(_753_), .C(_822_), .Y(_823_) );
AOI21X1 AOI21X1_146 ( .gnd(gnd), .vdd(vdd), .A(_823_), .B(_821_), .C(_786_), .Y(_824_) );
NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(_787_), .B(_822_), .Y(_825_) );
AOI21X1 AOI21X1_147 ( .gnd(gnd), .vdd(vdd), .A(_817_), .B(_819_), .C(_787_), .Y(_826_) );
INVX1 INVX1_631 ( .gnd(gnd), .vdd(vdd), .A(_826_), .Y(_827_) );
AOI21X1 AOI21X1_148 ( .gnd(gnd), .vdd(vdd), .A(_827_), .B(_825_), .C(_785_), .Y(_828_) );
OAI21X1 OAI21X1_815 ( .gnd(gnd), .vdd(vdd), .A(_824_), .B(_828_), .C(_784_), .Y(_829_) );
NAND3X1 NAND3X1_230 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_825_), .C(_827_), .Y(_830_) );
NAND3X1 NAND3X1_231 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_821_), .C(_823_), .Y(_831_) );
NAND3X1 NAND3X1_232 ( .gnd(gnd), .vdd(vdd), .A(_783_), .B(_831_), .C(_830_), .Y(_832_) );
AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_829_), .B(_832_), .Y(_833_) );
OAI21X1 OAI21X1_816 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_776_), .C(_833_), .Y(_834_) );
INVX1 INVX1_632 ( .gnd(gnd), .vdd(vdd), .A(_834_), .Y(_835_) );
NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_507_), .B(_777_), .Y(_836_) );
AOI21X1 AOI21X1_149 ( .gnd(gnd), .vdd(vdd), .A(_241_), .B(_836_), .C(_782_), .Y(_837_) );
INVX1 INVX1_633 ( .gnd(gnd), .vdd(vdd), .A(_837_), .Y(_838_) );
OAI21X1 OAI21X1_817 ( .gnd(gnd), .vdd(vdd), .A(_833_), .B(_838_), .C(round_ctr_inc_bF_buf9), .Y(_839_) );
INVX1 INVX1_634 ( .gnd(gnd), .vdd(vdd), .A(_3667__144_), .Y(_840_) );
OAI21X1 OAI21X1_818 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_840_), .Y(_841_) );
AOI22X1 AOI22X1_648 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf7), .B(_841_), .C(a_reg_16_), .D(_113__bF_buf0), .Y(_842_) );
OAI21X1 OAI21X1_819 ( .gnd(gnd), .vdd(vdd), .A(_835_), .B(_839_), .C(_842_), .Y(_5__16_) );
INVX2 INVX2_35 ( .gnd(gnd), .vdd(vdd), .A(a_reg_17_), .Y(_843_) );
INVX1 INVX1_635 ( .gnd(gnd), .vdd(vdd), .A(_832_), .Y(_844_) );
OAI21X1 OAI21X1_820 ( .gnd(gnd), .vdd(vdd), .A(_816_), .B(_801_), .C(_815_), .Y(_845_) );
INVX2 INVX2_36 ( .gnd(gnd), .vdd(vdd), .A(b_reg_17_), .Y(_846_) );
INVX2 INVX2_37 ( .gnd(gnd), .vdd(vdd), .A(c_reg_17_), .Y(_847_) );
NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_846_), .Y(_848_) );
AOI21X1 AOI21X1_150 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(d_reg_17_), .C(_848_), .Y(_849_) );
OAI21X1 OAI21X1_821 ( .gnd(gnd), .vdd(vdd), .A(c_reg_17_), .B(b_reg_17_), .C(d_reg_17_), .Y(_850_) );
OAI21X1 OAI21X1_822 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_846_), .C(_850_), .Y(_851_) );
NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_851_), .B(_3451__bF_buf0), .Y(_852_) );
INVX1 INVX1_636 ( .gnd(gnd), .vdd(vdd), .A(d_reg_17_), .Y(_853_) );
NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(c_reg_17_), .B(b_reg_17_), .Y(_854_) );
NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(d_reg_17_), .B(_848_), .Y(_855_) );
AOI22X1 AOI22X1_649 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_854_), .C(_851_), .D(_855_), .Y(_856_) );
AOI21X1 AOI21X1_151 ( .gnd(gnd), .vdd(vdd), .A(_856_), .B(_3405__bF_buf1), .C(_3447__bF_buf1), .Y(_857_) );
AOI22X1 AOI22X1_650 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf0), .B(_849_), .C(_852_), .D(_857_), .Y(_858_) );
INVX1 INVX1_637 ( .gnd(gnd), .vdd(vdd), .A(_805_), .Y(_859_) );
AOI21X1 AOI21X1_152 ( .gnd(gnd), .vdd(vdd), .A(_808_), .B(w_16_), .C(_859_), .Y(_860_) );
INVX1 INVX1_638 ( .gnd(gnd), .vdd(vdd), .A(_860_), .Y(_861_) );
INVX1 INVX1_639 ( .gnd(gnd), .vdd(vdd), .A(w_17_), .Y(_862_) );
NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(a_reg_12_), .B(e_reg_17_), .Y(_863_) );
INVX2 INVX2_38 ( .gnd(gnd), .vdd(vdd), .A(_863_), .Y(_864_) );
NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(a_reg_12_), .B(e_reg_17_), .Y(_865_) );
NOR3X1 NOR3X1_74 ( .gnd(gnd), .vdd(vdd), .A(_862_), .B(_865_), .C(_864_), .Y(_866_) );
INVX1 INVX1_640 ( .gnd(gnd), .vdd(vdd), .A(_866_), .Y(_867_) );
OAI21X1 OAI21X1_823 ( .gnd(gnd), .vdd(vdd), .A(_865_), .B(_864_), .C(_862_), .Y(_868_) );
NAND3X1 NAND3X1_233 ( .gnd(gnd), .vdd(vdd), .A(_868_), .B(_861_), .C(_867_), .Y(_869_) );
INVX1 INVX1_641 ( .gnd(gnd), .vdd(vdd), .A(_868_), .Y(_870_) );
OAI21X1 OAI21X1_824 ( .gnd(gnd), .vdd(vdd), .A(_866_), .B(_870_), .C(_860_), .Y(_871_) );
AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_869_), .B(_871_), .Y(_872_) );
NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_858_), .Y(_873_) );
AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_872_), .Y(_874_) );
OAI21X1 OAI21X1_825 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_874_), .C(_845_), .Y(_875_) );
INVX1 INVX1_642 ( .gnd(gnd), .vdd(vdd), .A(_815_), .Y(_876_) );
AOI21X1 AOI21X1_153 ( .gnd(gnd), .vdd(vdd), .A(_818_), .B(_812_), .C(_876_), .Y(_877_) );
OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_858_), .B(_872_), .Y(_878_) );
NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(_872_), .B(_858_), .Y(_879_) );
NAND3X1 NAND3X1_234 ( .gnd(gnd), .vdd(vdd), .A(_877_), .B(_879_), .C(_878_), .Y(_880_) );
NAND3X1 NAND3X1_235 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf0), .B(_880_), .C(_875_), .Y(_881_) );
NAND3X1 NAND3X1_236 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_845_), .C(_878_), .Y(_882_) );
OAI21X1 OAI21X1_826 ( .gnd(gnd), .vdd(vdd), .A(_873_), .B(_874_), .C(_877_), .Y(_883_) );
NAND3X1 NAND3X1_237 ( .gnd(gnd), .vdd(vdd), .A(_3473_), .B(_882_), .C(_883_), .Y(_884_) );
NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_884_), .Y(_885_) );
NAND3X1 NAND3X1_238 ( .gnd(gnd), .vdd(vdd), .A(_825_), .B(_830_), .C(_885_), .Y(_886_) );
OAI21X1 OAI21X1_827 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_826_), .C(_825_), .Y(_887_) );
NAND3X1 NAND3X1_239 ( .gnd(gnd), .vdd(vdd), .A(_881_), .B(_887_), .C(_884_), .Y(_888_) );
AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_888_), .Y(_889_) );
OAI21X1 OAI21X1_828 ( .gnd(gnd), .vdd(vdd), .A(_844_), .B(_835_), .C(_889_), .Y(_890_) );
NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_886_), .Y(_891_) );
NAND3X1 NAND3X1_240 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_891_), .C(_834_), .Y(_892_) );
AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_892_), .B(round_ctr_inc_bF_buf8), .Y(_893_) );
INVX2 INVX2_39 ( .gnd(gnd), .vdd(vdd), .A(_3667__145_), .Y(_894_) );
NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_3432__bF_buf9), .Y(_895_) );
AOI22X1 AOI22X1_651 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf6), .B(_895_), .C(_890_), .D(_893_), .Y(_896_) );
OAI21X1 OAI21X1_829 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_3387__bF_buf2), .C(_896_), .Y(_5__17_) );
NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(_888_), .B(_832_), .Y(_897_) );
NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_886_), .B(_897_), .Y(_898_) );
OAI21X1 OAI21X1_830 ( .gnd(gnd), .vdd(vdd), .A(_891_), .B(_834_), .C(_898_), .Y(_899_) );
AOI21X1 AOI21X1_154 ( .gnd(gnd), .vdd(vdd), .A(_878_), .B(_879_), .C(_845_), .Y(_900_) );
OAI21X1 OAI21X1_831 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf3), .B(_900_), .C(_882_), .Y(_901_) );
AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_879_), .B(_869_), .Y(_902_) );
INVX2 INVX2_40 ( .gnd(gnd), .vdd(vdd), .A(d_reg_18_), .Y(_903_) );
XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(c_reg_18_), .B(b_reg_18_), .Y(_904_) );
NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_904_), .Y(_905_) );
AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_904_), .B(_903_), .Y(_906_) );
OAI21X1 OAI21X1_832 ( .gnd(gnd), .vdd(vdd), .A(_905_), .B(_906_), .C(_3474__bF_buf2), .Y(_907_) );
INVX1 INVX1_643 ( .gnd(gnd), .vdd(vdd), .A(c_reg_18_), .Y(_908_) );
INVX2 INVX2_41 ( .gnd(gnd), .vdd(vdd), .A(b_reg_18_), .Y(_909_) );
OAI21X1 OAI21X1_833 ( .gnd(gnd), .vdd(vdd), .A(_908_), .B(_909_), .C(_903_), .Y(_910_) );
OAI21X1 OAI21X1_834 ( .gnd(gnd), .vdd(vdd), .A(c_reg_18_), .B(b_reg_18_), .C(_910_), .Y(_911_) );
NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(_911_), .B(_3405__bF_buf0), .Y(_912_) );
OAI21X1 OAI21X1_835 ( .gnd(gnd), .vdd(vdd), .A(c_reg_18_), .B(_909_), .C(_910_), .Y(_913_) );
NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf1), .B(_913_), .Y(_914_) );
NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_914_), .B(_912_), .Y(_915_) );
NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_907_), .B(_915_), .Y(_916_) );
NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_866_), .Y(_917_) );
INVX1 INVX1_644 ( .gnd(gnd), .vdd(vdd), .A(a_reg_13_), .Y(_918_) );
INVX1 INVX1_645 ( .gnd(gnd), .vdd(vdd), .A(e_reg_18_), .Y(_919_) );
NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_918_), .B(_919_), .Y(_920_) );
NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(a_reg_13_), .B(e_reg_18_), .Y(_921_) );
NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_921_), .B(_920_), .Y(_922_) );
AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(w_18_), .Y(_923_) );
NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(w_18_), .B(_922_), .Y(_924_) );
OAI21X1 OAI21X1_836 ( .gnd(gnd), .vdd(vdd), .A(_924_), .B(_923_), .C(_917_), .Y(_925_) );
INVX1 INVX1_646 ( .gnd(gnd), .vdd(vdd), .A(w_18_), .Y(_926_) );
XNOR2X1 XNOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(_922_), .B(_926_), .Y(_927_) );
OAI21X1 OAI21X1_837 ( .gnd(gnd), .vdd(vdd), .A(_864_), .B(_866_), .C(_927_), .Y(_928_) );
NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(_925_), .B(_928_), .Y(_929_) );
XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_916_), .Y(_930_) );
NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_902_), .B(_930_), .Y(_931_) );
INVX1 INVX1_647 ( .gnd(gnd), .vdd(vdd), .A(_869_), .Y(_932_) );
XNOR2X1 XNOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_916_), .Y(_933_) );
OAI21X1 OAI21X1_838 ( .gnd(gnd), .vdd(vdd), .A(_932_), .B(_874_), .C(_933_), .Y(_934_) );
NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_934_), .Y(_935_) );
NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_935_), .Y(_936_) );
OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_901_), .Y(_937_) );
NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_936_), .B(_937_), .Y(_938_) );
AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_899_), .B(_938_), .Y(_939_) );
OAI21X1 OAI21X1_839 ( .gnd(gnd), .vdd(vdd), .A(_938_), .B(_899_), .C(round_ctr_inc_bF_buf7), .Y(_940_) );
INVX1 INVX1_648 ( .gnd(gnd), .vdd(vdd), .A(_3667__146_), .Y(_941_) );
OAI21X1 OAI21X1_840 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_941_), .Y(_942_) );
AOI22X1 AOI22X1_652 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf5), .B(_942_), .C(a_reg_18_), .D(_113__bF_buf4), .Y(_943_) );
OAI21X1 OAI21X1_841 ( .gnd(gnd), .vdd(vdd), .A(_939_), .B(_940_), .C(_943_), .Y(_5__18_) );
NAND3X1 NAND3X1_241 ( .gnd(gnd), .vdd(vdd), .A(_931_), .B(_934_), .C(_901_), .Y(_944_) );
INVX1 INVX1_649 ( .gnd(gnd), .vdd(vdd), .A(_944_), .Y(_945_) );
NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(_945_), .B(_939_), .Y(_946_) );
INVX1 INVX1_650 ( .gnd(gnd), .vdd(vdd), .A(_916_), .Y(_947_) );
OAI21X1 OAI21X1_842 ( .gnd(gnd), .vdd(vdd), .A(_929_), .B(_947_), .C(_928_), .Y(_948_) );
INVX2 INVX2_42 ( .gnd(gnd), .vdd(vdd), .A(d_reg_19_), .Y(_949_) );
XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(c_reg_19_), .B(b_reg_19_), .Y(_950_) );
NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_950_), .Y(_951_) );
AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(_950_), .B(_949_), .Y(_952_) );
OAI21X1 OAI21X1_843 ( .gnd(gnd), .vdd(vdd), .A(_951_), .B(_952_), .C(_3474__bF_buf1), .Y(_953_) );
INVX1 INVX1_651 ( .gnd(gnd), .vdd(vdd), .A(c_reg_19_), .Y(_954_) );
INVX2 INVX2_43 ( .gnd(gnd), .vdd(vdd), .A(b_reg_19_), .Y(_955_) );
OAI21X1 OAI21X1_844 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_955_), .C(_949_), .Y(_956_) );
OAI21X1 OAI21X1_845 ( .gnd(gnd), .vdd(vdd), .A(c_reg_19_), .B(b_reg_19_), .C(_956_), .Y(_957_) );
NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_957_), .B(_3405__bF_buf5), .Y(_958_) );
OAI21X1 OAI21X1_846 ( .gnd(gnd), .vdd(vdd), .A(c_reg_19_), .B(_955_), .C(_956_), .Y(_959_) );
NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf0), .B(_959_), .Y(_960_) );
NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_960_), .B(_958_), .Y(_961_) );
NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_953_), .B(_961_), .Y(_962_) );
INVX1 INVX1_652 ( .gnd(gnd), .vdd(vdd), .A(_920_), .Y(_963_) );
OAI21X1 OAI21X1_847 ( .gnd(gnd), .vdd(vdd), .A(_926_), .B(_921_), .C(_963_), .Y(_964_) );
INVX1 INVX1_653 ( .gnd(gnd), .vdd(vdd), .A(_964_), .Y(_965_) );
NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(a_reg_14_), .B(e_reg_19_), .Y(_966_) );
INVX1 INVX1_654 ( .gnd(gnd), .vdd(vdd), .A(_966_), .Y(_967_) );
NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(a_reg_14_), .B(e_reg_19_), .Y(_968_) );
NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_967_), .Y(_969_) );
NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(w_19_), .B(_969_), .Y(_970_) );
INVX1 INVX1_655 ( .gnd(gnd), .vdd(vdd), .A(w_19_), .Y(_971_) );
OAI21X1 OAI21X1_848 ( .gnd(gnd), .vdd(vdd), .A(_968_), .B(_967_), .C(_971_), .Y(_972_) );
NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_970_), .Y(_973_) );
NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_965_), .B(_973_), .Y(_974_) );
NAND3X1 NAND3X1_242 ( .gnd(gnd), .vdd(vdd), .A(_972_), .B(_964_), .C(_970_), .Y(_975_) );
NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_975_), .B(_974_), .Y(_976_) );
XNOR2X1 XNOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_962_), .Y(_977_) );
NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(_948_), .B(_977_), .Y(_978_) );
INVX1 INVX1_656 ( .gnd(gnd), .vdd(vdd), .A(_928_), .Y(_979_) );
AOI21X1 AOI21X1_155 ( .gnd(gnd), .vdd(vdd), .A(_916_), .B(_925_), .C(_979_), .Y(_980_) );
AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_974_), .B(_975_), .Y(_981_) );
NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_981_), .Y(_982_) );
INVX1 INVX1_657 ( .gnd(gnd), .vdd(vdd), .A(_962_), .Y(_983_) );
NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_983_), .Y(_984_) );
OAI21X1 OAI21X1_849 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_984_), .C(_980_), .Y(_985_) );
NAND3X1 NAND3X1_243 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_985_), .C(_978_), .Y(_986_) );
NOR3X1 NOR3X1_75 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_980_), .C(_984_), .Y(_987_) );
NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_983_), .Y(_988_) );
NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_981_), .Y(_989_) );
AOI21X1 AOI21X1_156 ( .gnd(gnd), .vdd(vdd), .A(_989_), .B(_988_), .C(_948_), .Y(_990_) );
OAI21X1 OAI21X1_850 ( .gnd(gnd), .vdd(vdd), .A(_990_), .B(_987_), .C(_786_), .Y(_991_) );
NAND3X1 NAND3X1_244 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_986_), .C(_991_), .Y(_992_) );
INVX1 INVX1_658 ( .gnd(gnd), .vdd(vdd), .A(_934_), .Y(_993_) );
OAI21X1 OAI21X1_851 ( .gnd(gnd), .vdd(vdd), .A(_982_), .B(_984_), .C(_948_), .Y(_994_) );
NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_980_), .B(_977_), .Y(_995_) );
NAND3X1 NAND3X1_245 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_994_), .C(_995_), .Y(_996_) );
NAND3X1 NAND3X1_246 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_985_), .C(_978_), .Y(_997_) );
NAND3X1 NAND3X1_247 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_993_), .C(_997_), .Y(_998_) );
NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(_998_), .B(_992_), .Y(_999_) );
INVX1 INVX1_659 ( .gnd(gnd), .vdd(vdd), .A(_999_), .Y(_1000_) );
AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(_946_), .B(_1000_), .Y(_1001_) );
OAI21X1 OAI21X1_852 ( .gnd(gnd), .vdd(vdd), .A(_1000_), .B(_946_), .C(round_ctr_inc_bF_buf6), .Y(_1002_) );
INVX1 INVX1_660 ( .gnd(gnd), .vdd(vdd), .A(_3667__147_), .Y(_1003_) );
NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .B(_3432__bF_buf8), .Y(_1004_) );
AOI22X1 AOI22X1_653 ( .gnd(gnd), .vdd(vdd), .A(_1004_), .B(_3433__bF_buf4), .C(a_reg_19_), .D(_113__bF_buf3), .Y(_1005_) );
OAI21X1 OAI21X1_853 ( .gnd(gnd), .vdd(vdd), .A(_1001_), .B(_1002_), .C(_1005_), .Y(_5__19_) );
NAND3X1 NAND3X1_248 ( .gnd(gnd), .vdd(vdd), .A(_934_), .B(_997_), .C(_996_), .Y(_1006_) );
NAND3X1 NAND3X1_249 ( .gnd(gnd), .vdd(vdd), .A(_993_), .B(_986_), .C(_991_), .Y(_1007_) );
NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_944_), .B(_1007_), .Y(_1008_) );
NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_1006_), .B(_1008_), .Y(_1009_) );
AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(_935_), .B(_901_), .Y(_1010_) );
NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_901_), .B(_935_), .Y(_1011_) );
AOI21X1 AOI21X1_157 ( .gnd(gnd), .vdd(vdd), .A(_996_), .B(_997_), .C(_993_), .Y(_1012_) );
AOI21X1 AOI21X1_158 ( .gnd(gnd), .vdd(vdd), .A(_991_), .B(_986_), .C(_934_), .Y(_1013_) );
OAI22X1 OAI22X1_55 ( .gnd(gnd), .vdd(vdd), .A(_1011_), .B(_1010_), .C(_1012_), .D(_1013_), .Y(_1014_) );
OAI21X1 OAI21X1_854 ( .gnd(gnd), .vdd(vdd), .A(_898_), .B(_1014_), .C(_1009_), .Y(_1015_) );
INVX1 INVX1_661 ( .gnd(gnd), .vdd(vdd), .A(_1015_), .Y(_1016_) );
AOI22X1 AOI22X1_654 ( .gnd(gnd), .vdd(vdd), .A(_992_), .B(_998_), .C(_936_), .D(_937_), .Y(_1017_) );
NAND3X1 NAND3X1_250 ( .gnd(gnd), .vdd(vdd), .A(_833_), .B(_1017_), .C(_889_), .Y(_1018_) );
OAI21X1 OAI21X1_855 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_837_), .C(_1016_), .Y(_1019_) );
OAI21X1 OAI21X1_856 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_990_), .C(_978_), .Y(_1020_) );
OAI21X1 OAI21X1_857 ( .gnd(gnd), .vdd(vdd), .A(_976_), .B(_983_), .C(_975_), .Y(_1021_) );
INVX2 INVX2_44 ( .gnd(gnd), .vdd(vdd), .A(c_reg_20_), .Y(_1022_) );
INVX2 INVX2_45 ( .gnd(gnd), .vdd(vdd), .A(b_reg_20_), .Y(_1023_) );
INVX1 INVX1_662 ( .gnd(gnd), .vdd(vdd), .A(d_reg_20_), .Y(_1024_) );
OAI21X1 OAI21X1_858 ( .gnd(gnd), .vdd(vdd), .A(_1022_), .B(_1023_), .C(_1024_), .Y(_1025_) );
OAI21X1 OAI21X1_859 ( .gnd(gnd), .vdd(vdd), .A(c_reg_20_), .B(b_reg_20_), .C(_1025_), .Y(_1026_) );
OAI21X1 OAI21X1_860 ( .gnd(gnd), .vdd(vdd), .A(c_reg_20_), .B(_1023_), .C(_1025_), .Y(_1027_) );
NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf4), .B(_1027_), .Y(_1028_) );
XNOR2X1 XNOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(c_reg_20_), .B(b_reg_20_), .Y(_1029_) );
XNOR2X1 XNOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1029_), .B(d_reg_20_), .Y(_1030_) );
AOI21X1 AOI21X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_3474__bF_buf0), .C(_1028_), .Y(_1031_) );
OAI21X1 OAI21X1_861 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf4), .B(_1026_), .C(_1031_), .Y(_1032_) );
OAI21X1 OAI21X1_862 ( .gnd(gnd), .vdd(vdd), .A(_971_), .B(_968_), .C(_966_), .Y(_1033_) );
INVX1 INVX1_663 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .Y(_1034_) );
NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(a_reg_15_), .B(e_reg_20_), .Y(_1035_) );
INVX1 INVX1_664 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .Y(_1036_) );
NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(a_reg_15_), .B(e_reg_20_), .Y(_1037_) );
NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .B(_1036_), .Y(_1038_) );
NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(w_20_), .B(_1038_), .Y(_1039_) );
INVX1 INVX1_665 ( .gnd(gnd), .vdd(vdd), .A(w_20_), .Y(_1040_) );
OAI21X1 OAI21X1_863 ( .gnd(gnd), .vdd(vdd), .A(_1037_), .B(_1036_), .C(_1040_), .Y(_1041_) );
NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_1041_), .B(_1039_), .Y(_1042_) );
NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_1034_), .B(_1042_), .Y(_1043_) );
NAND3X1 NAND3X1_251 ( .gnd(gnd), .vdd(vdd), .A(_1033_), .B(_1041_), .C(_1039_), .Y(_1044_) );
AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_1043_), .B(_1044_), .Y(_1045_) );
NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1032_), .Y(_1046_) );
OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf3), .B(_1026_), .Y(_1047_) );
OAI21X1 OAI21X1_864 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf3), .B(_1027_), .C(_1047_), .Y(_1048_) );
AOI21X1 AOI21X1_160 ( .gnd(gnd), .vdd(vdd), .A(_1030_), .B(_3474__bF_buf4), .C(_1048_), .Y(_1049_) );
NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .B(_1043_), .Y(_1050_) );
NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1049_), .Y(_1051_) );
OAI21X1 OAI21X1_865 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_1046_), .C(_1021_), .Y(_1052_) );
INVX1 INVX1_666 ( .gnd(gnd), .vdd(vdd), .A(_975_), .Y(_1053_) );
AOI21X1 AOI21X1_161 ( .gnd(gnd), .vdd(vdd), .A(_962_), .B(_974_), .C(_1053_), .Y(_1054_) );
NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1049_), .Y(_1055_) );
NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_1045_), .B(_1032_), .Y(_1056_) );
NAND3X1 NAND3X1_252 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1054_), .C(_1056_), .Y(_1057_) );
AOI21X1 AOI21X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1052_), .B(_1057_), .C(_786_), .Y(_1058_) );
NAND3X1 NAND3X1_253 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1056_), .C(_1021_), .Y(_1059_) );
OAI21X1 OAI21X1_866 ( .gnd(gnd), .vdd(vdd), .A(_1051_), .B(_1046_), .C(_1054_), .Y(_1060_) );
AOI21X1 AOI21X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1059_), .B(_1060_), .C(_785_), .Y(_1061_) );
OAI21X1 OAI21X1_867 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1061_), .C(_1020_), .Y(_1062_) );
AOI21X1 AOI21X1_164 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_985_), .C(_987_), .Y(_1063_) );
NAND3X1 NAND3X1_254 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_1060_), .C(_1059_), .Y(_1064_) );
NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_1055_), .B(_1056_), .Y(_1065_) );
NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1054_), .B(_1065_), .Y(_1066_) );
AOI21X1 AOI21X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1056_), .B(_1055_), .C(_1021_), .Y(_1067_) );
OAI21X1 OAI21X1_868 ( .gnd(gnd), .vdd(vdd), .A(_1067_), .B(_1066_), .C(_786_), .Y(_1068_) );
NAND3X1 NAND3X1_255 ( .gnd(gnd), .vdd(vdd), .A(_1063_), .B(_1064_), .C(_1068_), .Y(_1069_) );
NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_1062_), .B(_1069_), .Y(_1070_) );
XNOR2X1 XNOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1070_), .Y(_1071_) );
INVX1 INVX1_667 ( .gnd(gnd), .vdd(vdd), .A(_3667__148_), .Y(_1072_) );
NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_3432__bF_buf7), .Y(_1073_) );
AOI22X1 AOI22X1_655 ( .gnd(gnd), .vdd(vdd), .A(_1073_), .B(_3433__bF_buf3), .C(a_reg_20_), .D(_113__bF_buf2), .Y(_1074_) );
OAI21X1 OAI21X1_869 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_1071_), .C(_1074_), .Y(_5__20_) );
AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1070_), .Y(_1075_) );
NOR3X1 NOR3X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1061_), .C(_1063_), .Y(_1076_) );
INVX1 INVX1_668 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .Y(_1077_) );
AOI21X1 AOI21X1_166 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_1060_), .C(_1066_), .Y(_1078_) );
OAI21X1 OAI21X1_870 ( .gnd(gnd), .vdd(vdd), .A(_1050_), .B(_1049_), .C(_1044_), .Y(_1079_) );
XNOR2X1 XNOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(c_reg_21_), .B(b_reg_21_), .Y(_1080_) );
XNOR2X1 XNOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1080_), .B(d_reg_21_), .Y(_1081_) );
INVX1 INVX1_669 ( .gnd(gnd), .vdd(vdd), .A(c_reg_21_), .Y(_1082_) );
INVX2 INVX2_46 ( .gnd(gnd), .vdd(vdd), .A(b_reg_21_), .Y(_1083_) );
INVX1 INVX1_670 ( .gnd(gnd), .vdd(vdd), .A(d_reg_21_), .Y(_1084_) );
OAI21X1 OAI21X1_871 ( .gnd(gnd), .vdd(vdd), .A(_1082_), .B(_1083_), .C(_1084_), .Y(_1085_) );
OAI21X1 OAI21X1_872 ( .gnd(gnd), .vdd(vdd), .A(c_reg_21_), .B(b_reg_21_), .C(_1085_), .Y(_1086_) );
OAI21X1 OAI21X1_873 ( .gnd(gnd), .vdd(vdd), .A(c_reg_21_), .B(_1083_), .C(_1085_), .Y(_1087_) );
OAI22X1 OAI22X1_56 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf2), .B(_1087_), .C(_1086_), .D(_3405__bF_buf2), .Y(_1088_) );
AOI21X1 AOI21X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1081_), .B(_3474__bF_buf3), .C(_1088_), .Y(_1089_) );
INVX1 INVX1_671 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .Y(_1090_) );
NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(a_reg_16_), .B(e_reg_21_), .Y(_1091_) );
INVX1 INVX1_672 ( .gnd(gnd), .vdd(vdd), .A(_1091_), .Y(_1092_) );
NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(a_reg_16_), .B(e_reg_21_), .Y(_1093_) );
NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1092_), .Y(_1094_) );
NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(w_21_), .B(_1094_), .Y(_1095_) );
INVX1 INVX1_673 ( .gnd(gnd), .vdd(vdd), .A(w_21_), .Y(_1096_) );
OAI21X1 OAI21X1_874 ( .gnd(gnd), .vdd(vdd), .A(_1093_), .B(_1092_), .C(_1096_), .Y(_1097_) );
NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_1097_), .B(_1095_), .Y(_1098_) );
NAND3X1 NAND3X1_256 ( .gnd(gnd), .vdd(vdd), .A(_1035_), .B(_1039_), .C(_1098_), .Y(_1099_) );
OAI21X1 OAI21X1_875 ( .gnd(gnd), .vdd(vdd), .A(_1040_), .B(_1037_), .C(_1035_), .Y(_1100_) );
NAND3X1 NAND3X1_257 ( .gnd(gnd), .vdd(vdd), .A(_1100_), .B(_1097_), .C(_1095_), .Y(_1101_) );
AOI21X1 AOI21X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1099_), .B(_1101_), .C(_1090_), .Y(_1102_) );
NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .B(_1099_), .Y(_1103_) );
NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1103_), .Y(_1104_) );
OAI21X1 OAI21X1_876 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_1102_), .C(_1079_), .Y(_1105_) );
INVX1 INVX1_674 ( .gnd(gnd), .vdd(vdd), .A(_1044_), .Y(_1106_) );
AOI21X1 AOI21X1_169 ( .gnd(gnd), .vdd(vdd), .A(_1032_), .B(_1043_), .C(_1106_), .Y(_1107_) );
NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1103_), .Y(_1108_) );
OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(_1103_), .B(_1089_), .Y(_1109_) );
NAND3X1 NAND3X1_258 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_1109_), .C(_1107_), .Y(_1110_) );
AOI21X1 AOI21X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1110_), .B(_1105_), .C(_3472_), .Y(_1111_) );
NAND3X1 NAND3X1_259 ( .gnd(gnd), .vdd(vdd), .A(_1108_), .B(_1079_), .C(_1109_), .Y(_1112_) );
OAI21X1 OAI21X1_877 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_1102_), .C(_1107_), .Y(_1113_) );
AOI21X1 AOI21X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1112_), .B(_1113_), .C(_3437__bF_buf1), .Y(_1114_) );
NOR3X1 NOR3X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_1111_), .C(_1078_), .Y(_1115_) );
OAI21X1 OAI21X1_878 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_1111_), .C(_1078_), .Y(_1116_) );
INVX1 INVX1_675 ( .gnd(gnd), .vdd(vdd), .A(_1116_), .Y(_1117_) );
OAI21X1 OAI21X1_879 ( .gnd(gnd), .vdd(vdd), .A(_1115_), .B(_1117_), .C(_1077_), .Y(_1118_) );
NAND3X1 NAND3X1_260 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf0), .B(_1113_), .C(_1112_), .Y(_1119_) );
NOR3X1 NOR3X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1104_), .B(_1102_), .C(_1107_), .Y(_1120_) );
AOI21X1 AOI21X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1109_), .B(_1108_), .C(_1079_), .Y(_1121_) );
OAI21X1 OAI21X1_880 ( .gnd(gnd), .vdd(vdd), .A(_1121_), .B(_1120_), .C(_3472_), .Y(_1122_) );
AOI21X1 AOI21X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1122_), .B(_1119_), .C(_1078_), .Y(_1123_) );
OAI21X1 OAI21X1_881 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_1067_), .C(_1059_), .Y(_1124_) );
NOR3X1 NOR3X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_1111_), .C(_1124_), .Y(_1125_) );
OAI22X1 OAI22X1_57 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1125_), .C(_1076_), .D(_1075_), .Y(_1126_) );
OAI21X1 OAI21X1_882 ( .gnd(gnd), .vdd(vdd), .A(_1075_), .B(_1118_), .C(_1126_), .Y(_1127_) );
INVX1 INVX1_676 ( .gnd(gnd), .vdd(vdd), .A(_3667__149_), .Y(_1128_) );
NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_3432__bF_buf6), .Y(_1129_) );
AOI22X1 AOI22X1_656 ( .gnd(gnd), .vdd(vdd), .A(_1129_), .B(_3433__bF_buf2), .C(a_reg_21_), .D(_113__bF_buf1), .Y(_1130_) );
OAI21X1 OAI21X1_883 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_1127_), .C(_1130_), .Y(_5__21_) );
OAI21X1 OAI21X1_884 ( .gnd(gnd), .vdd(vdd), .A(_1114_), .B(_1111_), .C(_1124_), .Y(_1131_) );
NAND3X1 NAND3X1_261 ( .gnd(gnd), .vdd(vdd), .A(_1119_), .B(_1078_), .C(_1122_), .Y(_1132_) );
AOI22X1 AOI22X1_657 ( .gnd(gnd), .vdd(vdd), .A(_1132_), .B(_1131_), .C(_1062_), .D(_1069_), .Y(_1133_) );
AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(_1019_), .B(_1133_), .Y(_1134_) );
AOI21X1 AOI21X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1076_), .B(_1116_), .C(_1115_), .Y(_1135_) );
INVX1 INVX1_677 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .Y(_1136_) );
NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1136_), .B(_1134_), .Y(_1137_) );
OAI21X1 OAI21X1_885 ( .gnd(gnd), .vdd(vdd), .A(_3472_), .B(_1121_), .C(_1112_), .Y(_1138_) );
OAI21X1 OAI21X1_886 ( .gnd(gnd), .vdd(vdd), .A(_1089_), .B(_1103_), .C(_1101_), .Y(_1139_) );
INVX2 INVX2_47 ( .gnd(gnd), .vdd(vdd), .A(c_reg_22_), .Y(_1140_) );
INVX2 INVX2_48 ( .gnd(gnd), .vdd(vdd), .A(b_reg_22_), .Y(_1141_) );
INVX2 INVX2_49 ( .gnd(gnd), .vdd(vdd), .A(d_reg_22_), .Y(_1142_) );
OAI21X1 OAI21X1_887 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1141_), .C(_1142_), .Y(_1143_) );
OAI21X1 OAI21X1_888 ( .gnd(gnd), .vdd(vdd), .A(c_reg_22_), .B(b_reg_22_), .C(_1143_), .Y(_1144_) );
NAND3X1 NAND3X1_262 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1141_), .C(_1142_), .Y(_1145_) );
NAND3X1 NAND3X1_263 ( .gnd(gnd), .vdd(vdd), .A(c_reg_22_), .B(b_reg_22_), .C(d_reg_22_), .Y(_1146_) );
INVX1 INVX1_678 ( .gnd(gnd), .vdd(vdd), .A(_1146_), .Y(_1147_) );
OAI21X1 OAI21X1_889 ( .gnd(gnd), .vdd(vdd), .A(_1147_), .B(_1144_), .C(_1145_), .Y(_1148_) );
NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1144_), .B(_3405__bF_buf1), .Y(_1149_) );
OAI21X1 OAI21X1_890 ( .gnd(gnd), .vdd(vdd), .A(c_reg_22_), .B(_1141_), .C(_1143_), .Y(_1150_) );
NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_3411__bF_buf1), .B(_1150_), .Y(_1151_) );
NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1151_), .B(_1149_), .Y(_1152_) );
OAI21X1 OAI21X1_891 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf1), .B(_1148_), .C(_1152_), .Y(_1153_) );
OAI21X1 OAI21X1_892 ( .gnd(gnd), .vdd(vdd), .A(_1096_), .B(_1093_), .C(_1091_), .Y(_1154_) );
INVX1 INVX1_679 ( .gnd(gnd), .vdd(vdd), .A(_1154_), .Y(_1155_) );
INVX1 INVX1_680 ( .gnd(gnd), .vdd(vdd), .A(w_22_), .Y(_1156_) );
INVX1 INVX1_681 ( .gnd(gnd), .vdd(vdd), .A(e_reg_22_), .Y(_1157_) );
NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_843_), .B(_1157_), .Y(_1158_) );
NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(a_reg_17_), .B(e_reg_22_), .Y(_1159_) );
NOR3X1 NOR3X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1156_), .B(_1159_), .C(_1158_), .Y(_1160_) );
OAI21X1 OAI21X1_893 ( .gnd(gnd), .vdd(vdd), .A(_1159_), .B(_1158_), .C(_1156_), .Y(_1161_) );
INVX1 INVX1_682 ( .gnd(gnd), .vdd(vdd), .A(_1161_), .Y(_1162_) );
OAI21X1 OAI21X1_894 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .B(_1162_), .C(_1155_), .Y(_1163_) );
INVX1 INVX1_683 ( .gnd(gnd), .vdd(vdd), .A(_1160_), .Y(_1164_) );
NAND3X1 NAND3X1_264 ( .gnd(gnd), .vdd(vdd), .A(_1154_), .B(_1161_), .C(_1164_), .Y(_1165_) );
AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .B(_1163_), .Y(_1166_) );
NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1166_), .Y(_1167_) );
AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(_1166_), .B(_1153_), .Y(_1168_) );
OAI21X1 OAI21X1_895 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_1168_), .C(_1139_), .Y(_1169_) );
INVX1 INVX1_684 ( .gnd(gnd), .vdd(vdd), .A(_1101_), .Y(_1170_) );
AOI21X1 AOI21X1_175 ( .gnd(gnd), .vdd(vdd), .A(_1090_), .B(_1099_), .C(_1170_), .Y(_1171_) );
OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(_1166_), .B(_1153_), .Y(_1172_) );
NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1166_), .Y(_1173_) );
NAND3X1 NAND3X1_265 ( .gnd(gnd), .vdd(vdd), .A(_1173_), .B(_1171_), .C(_1172_), .Y(_1174_) );
AOI21X1 AOI21X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1169_), .B(_1174_), .C(_3406__bF_buf0), .Y(_1175_) );
NAND3X1 NAND3X1_266 ( .gnd(gnd), .vdd(vdd), .A(_1139_), .B(_1173_), .C(_1172_), .Y(_1176_) );
OAI21X1 OAI21X1_896 ( .gnd(gnd), .vdd(vdd), .A(_1167_), .B(_1168_), .C(_1171_), .Y(_1177_) );
AOI21X1 AOI21X1_177 ( .gnd(gnd), .vdd(vdd), .A(_1177_), .B(_1176_), .C(_3474__bF_buf2), .Y(_1178_) );
OAI21X1 OAI21X1_897 ( .gnd(gnd), .vdd(vdd), .A(_1175_), .B(_1178_), .C(_1138_), .Y(_1179_) );
AOI21X1 AOI21X1_178 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf3), .B(_1113_), .C(_1120_), .Y(_1180_) );
NAND3X1 NAND3X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3474__bF_buf1), .B(_1176_), .C(_1177_), .Y(_1181_) );
NAND3X1 NAND3X1_268 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf4), .B(_1174_), .C(_1169_), .Y(_1182_) );
NAND3X1 NAND3X1_269 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_1182_), .C(_1180_), .Y(_1183_) );
NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_1179_), .B(_1183_), .Y(_1184_) );
INVX1 INVX1_685 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .Y(_1185_) );
AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(_1137_), .B(_1185_), .Y(_1186_) );
OAI21X1 OAI21X1_898 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_1137_), .C(round_ctr_inc_bF_buf5), .Y(_1187_) );
INVX1 INVX1_686 ( .gnd(gnd), .vdd(vdd), .A(_3667__150_), .Y(_1188_) );
OAI21X1 OAI21X1_899 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1188_), .Y(_1189_) );
AOI22X1 AOI22X1_658 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf1), .B(_1189_), .C(a_reg_22_), .D(_113__bF_buf0), .Y(_1190_) );
OAI21X1 OAI21X1_900 ( .gnd(gnd), .vdd(vdd), .A(_1186_), .B(_1187_), .C(_1190_), .Y(_5__22_) );
NAND3X1 NAND3X1_270 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_1182_), .C(_1138_), .Y(_1191_) );
OAI21X1 OAI21X1_901 ( .gnd(gnd), .vdd(vdd), .A(_1185_), .B(_1137_), .C(_1191_), .Y(_1192_) );
NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_1176_), .B(_1181_), .Y(_1193_) );
INVX1 INVX1_687 ( .gnd(gnd), .vdd(vdd), .A(_1165_), .Y(_1194_) );
AOI21X1 AOI21X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1153_), .B(_1163_), .C(_1194_), .Y(_1195_) );
INVX1 INVX1_688 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .Y(_1196_) );
INVX2 INVX2_50 ( .gnd(gnd), .vdd(vdd), .A(b_reg_23_), .Y(_1197_) );
INVX2 INVX2_51 ( .gnd(gnd), .vdd(vdd), .A(c_reg_23_), .Y(_1198_) );
NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_1197_), .Y(_1199_) );
AOI21X1 AOI21X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(d_reg_23_), .C(_1199_), .Y(_1200_) );
NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf4), .B(_1200_), .Y(_1201_) );
OAI21X1 OAI21X1_902 ( .gnd(gnd), .vdd(vdd), .A(c_reg_23_), .B(b_reg_23_), .C(d_reg_23_), .Y(_1202_) );
OAI21X1 OAI21X1_903 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_1197_), .C(_1202_), .Y(_1203_) );
NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_1203_), .B(_3451__bF_buf4), .Y(_1204_) );
INVX1 INVX1_689 ( .gnd(gnd), .vdd(vdd), .A(d_reg_23_), .Y(_1205_) );
NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(c_reg_23_), .B(b_reg_23_), .Y(_1206_) );
NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(d_reg_23_), .B(_1199_), .Y(_1207_) );
AOI22X1 AOI22X1_659 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1206_), .C(_1203_), .D(_1207_), .Y(_1208_) );
AOI21X1 AOI21X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1208_), .B(_3405__bF_buf0), .C(_3447__bF_buf3), .Y(_1209_) );
NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_1204_), .B(_1209_), .Y(_1210_) );
NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(_1201_), .B(_1210_), .Y(_1211_) );
INVX1 INVX1_690 ( .gnd(gnd), .vdd(vdd), .A(_1158_), .Y(_1212_) );
OAI21X1 OAI21X1_904 ( .gnd(gnd), .vdd(vdd), .A(_1156_), .B(_1159_), .C(_1212_), .Y(_1213_) );
INVX1 INVX1_691 ( .gnd(gnd), .vdd(vdd), .A(a_reg_18_), .Y(_1214_) );
INVX1 INVX1_692 ( .gnd(gnd), .vdd(vdd), .A(e_reg_23_), .Y(_1215_) );
NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_1214_), .B(_1215_), .Y(_1216_) );
NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(a_reg_18_), .B(e_reg_23_), .Y(_1217_) );
NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_1217_), .B(_1216_), .Y(_1218_) );
NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(w_23_), .B(_1218_), .Y(_1219_) );
INVX1 INVX1_693 ( .gnd(gnd), .vdd(vdd), .A(w_23_), .Y(_1220_) );
OAI21X1 OAI21X1_905 ( .gnd(gnd), .vdd(vdd), .A(_1217_), .B(_1216_), .C(_1220_), .Y(_1221_) );
NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_1221_), .B(_1219_), .Y(_1222_) );
XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_1213_), .Y(_1223_) );
NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1211_), .Y(_1224_) );
AOI22X1 AOI22X1_660 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf2), .B(_1200_), .C(_1204_), .D(_1209_), .Y(_1225_) );
XNOR2X1 XNOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1222_), .B(_1213_), .Y(_1226_) );
NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_1226_), .Y(_1227_) );
AOI21X1 AOI21X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1227_), .C(_1196_), .Y(_1228_) );
NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_1225_), .B(_1226_), .Y(_1229_) );
NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_1223_), .B(_1211_), .Y(_1230_) );
NOR3X1 NOR3X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1195_), .B(_1229_), .C(_1230_), .Y(_1231_) );
OAI21X1 OAI21X1_906 ( .gnd(gnd), .vdd(vdd), .A(_1228_), .B(_1231_), .C(_3391_), .Y(_1232_) );
OAI21X1 OAI21X1_907 ( .gnd(gnd), .vdd(vdd), .A(_1229_), .B(_1230_), .C(_1195_), .Y(_1233_) );
NAND3X1 NAND3X1_271 ( .gnd(gnd), .vdd(vdd), .A(_1224_), .B(_1227_), .C(_1196_), .Y(_1234_) );
NAND3X1 NAND3X1_272 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_1234_), .C(_1233_), .Y(_1235_) );
NAND3X1 NAND3X1_273 ( .gnd(gnd), .vdd(vdd), .A(_1235_), .B(_1232_), .C(_1193_), .Y(_1236_) );
AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(_1181_), .B(_1176_), .Y(_1237_) );
AOI21X1 AOI21X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1233_), .B(_1234_), .C(_3392_), .Y(_1238_) );
NOR3X1 NOR3X1_82 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .B(_1228_), .C(_1231_), .Y(_1239_) );
OAI21X1 OAI21X1_908 ( .gnd(gnd), .vdd(vdd), .A(_1238_), .B(_1239_), .C(_1237_), .Y(_1240_) );
AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .B(_1236_), .Y(_1241_) );
AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(_1192_), .B(_1241_), .Y(_1242_) );
OAI21X1 OAI21X1_909 ( .gnd(gnd), .vdd(vdd), .A(_1241_), .B(_1192_), .C(round_ctr_inc_bF_buf4), .Y(_1243_) );
INVX1 INVX1_694 ( .gnd(gnd), .vdd(vdd), .A(_3667__151_), .Y(_1244_) );
NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_3432__bF_buf5), .Y(_1245_) );
AOI22X1 AOI22X1_661 ( .gnd(gnd), .vdd(vdd), .A(_1245_), .B(_3433__bF_buf0), .C(a_reg_23_), .D(_113__bF_buf4), .Y(_1246_) );
OAI21X1 OAI21X1_910 ( .gnd(gnd), .vdd(vdd), .A(_1242_), .B(_1243_), .C(_1246_), .Y(_5__23_) );
INVX1 INVX1_695 ( .gnd(gnd), .vdd(vdd), .A(a_reg_24_), .Y(_1247_) );
NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_832_), .B(_829_), .Y(_1248_) );
NOR3X1 NOR3X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1248_), .B(_891_), .C(_1014_), .Y(_1249_) );
AOI21X1 AOI21X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1068_), .B(_1064_), .C(_1063_), .Y(_1250_) );
NOR3X1 NOR3X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1058_), .B(_1061_), .C(_1020_), .Y(_1251_) );
OAI22X1 OAI22X1_58 ( .gnd(gnd), .vdd(vdd), .A(_1123_), .B(_1125_), .C(_1250_), .D(_1251_), .Y(_1252_) );
NAND3X1 NAND3X1_274 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .B(_1240_), .C(_1184_), .Y(_1253_) );
NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_1252_), .B(_1253_), .Y(_1254_) );
NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1249_), .Y(_1255_) );
INVX1 INVX1_696 ( .gnd(gnd), .vdd(vdd), .A(_1191_), .Y(_1256_) );
INVX1 INVX1_697 ( .gnd(gnd), .vdd(vdd), .A(_1236_), .Y(_1257_) );
AOI21X1 AOI21X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1240_), .B(_1256_), .C(_1257_), .Y(_1258_) );
OAI21X1 OAI21X1_911 ( .gnd(gnd), .vdd(vdd), .A(_1135_), .B(_1253_), .C(_1258_), .Y(_1259_) );
AOI21X1 AOI21X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1254_), .B(_1015_), .C(_1259_), .Y(_1260_) );
OAI21X1 OAI21X1_912 ( .gnd(gnd), .vdd(vdd), .A(_1255_), .B(_837_), .C(_1260_), .Y(_1261_) );
OAI21X1 OAI21X1_913 ( .gnd(gnd), .vdd(vdd), .A(_3391_), .B(_1228_), .C(_1234_), .Y(_1262_) );
INVX1 INVX1_698 ( .gnd(gnd), .vdd(vdd), .A(_1262_), .Y(_1263_) );
INVX1 INVX1_699 ( .gnd(gnd), .vdd(vdd), .A(_1213_), .Y(_1264_) );
OAI21X1 OAI21X1_914 ( .gnd(gnd), .vdd(vdd), .A(_1264_), .B(_1222_), .C(_1227_), .Y(_1265_) );
INVX2 INVX2_52 ( .gnd(gnd), .vdd(vdd), .A(b_reg_24_), .Y(_1266_) );
INVX1 INVX1_700 ( .gnd(gnd), .vdd(vdd), .A(c_reg_24_), .Y(_1267_) );
INVX2 INVX2_53 ( .gnd(gnd), .vdd(vdd), .A(d_reg_24_), .Y(_1268_) );
OAI21X1 OAI21X1_915 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1266_), .C(_1268_), .Y(_1269_) );
OAI21X1 OAI21X1_916 ( .gnd(gnd), .vdd(vdd), .A(c_reg_24_), .B(_1266_), .C(_1269_), .Y(_1270_) );
NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf1), .B(_1270_), .Y(_1271_) );
OAI21X1 OAI21X1_917 ( .gnd(gnd), .vdd(vdd), .A(c_reg_24_), .B(b_reg_24_), .C(_1269_), .Y(_1272_) );
XNOR2X1 XNOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(c_reg_24_), .B(b_reg_24_), .Y(_1273_) );
XNOR2X1 XNOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1273_), .B(_1268_), .Y(_1274_) );
OAI22X1 OAI22X1_59 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf5), .B(_1272_), .C(_3406__bF_buf3), .D(_1274_), .Y(_1275_) );
OAI21X1 OAI21X1_918 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf0), .B(_1275_), .C(_1271_), .Y(_1276_) );
INVX1 INVX1_701 ( .gnd(gnd), .vdd(vdd), .A(_1216_), .Y(_1277_) );
OAI21X1 OAI21X1_919 ( .gnd(gnd), .vdd(vdd), .A(_1220_), .B(_1217_), .C(_1277_), .Y(_1278_) );
INVX1 INVX1_702 ( .gnd(gnd), .vdd(vdd), .A(a_reg_19_), .Y(_1279_) );
INVX1 INVX1_703 ( .gnd(gnd), .vdd(vdd), .A(e_reg_24_), .Y(_1280_) );
NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_1279_), .B(_1280_), .Y(_1281_) );
NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(a_reg_19_), .B(e_reg_24_), .Y(_1282_) );
NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_1282_), .B(_1281_), .Y(_1283_) );
XNOR2X1 XNOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(w_24_), .Y(_1284_) );
XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .B(_1278_), .Y(_1285_) );
XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_1285_), .B(_1276_), .Y(_1286_) );
NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_1265_), .B(_1286_), .Y(_1287_) );
OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1265_), .Y(_1288_) );
NAND3X1 NAND3X1_275 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf3), .B(_1287_), .C(_1288_), .Y(_1289_) );
XNOR2X1 XNOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1286_), .B(_1265_), .Y(_1290_) );
OAI21X1 OAI21X1_920 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3437__bF_buf2), .C(_1290_), .Y(_1291_) );
AOI21X1 AOI21X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1291_), .B(_1289_), .C(_1263_), .Y(_1292_) );
INVX1 INVX1_704 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .Y(_1293_) );
NAND3X1 NAND3X1_276 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(_1289_), .C(_1291_), .Y(_1294_) );
NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .B(_1293_), .Y(_1295_) );
AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1295_), .Y(_1296_) );
NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_1296_), .Y(_1297_) );
OAI21X1 OAI21X1_921 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1295_), .C(_1297_), .Y(_1298_) );
OAI21X1 OAI21X1_922 ( .gnd(gnd), .vdd(vdd), .A(_3667__152_), .B(_3432__bF_buf4), .C(_3433__bF_buf11), .Y(_1299_) );
AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(_1298_), .B(_1299_), .Y(_1300_) );
OAI21X1 OAI21X1_923 ( .gnd(gnd), .vdd(vdd), .A(_1247_), .B(_3387__bF_buf1), .C(_1300_), .Y(_5__24_) );
NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_1289_), .B(_1291_), .Y(_1301_) );
NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_1263_), .B(_1301_), .Y(_1302_) );
OAI21X1 OAI21X1_924 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf4), .B(_1290_), .C(_1287_), .Y(_1303_) );
INVX1 INVX1_705 ( .gnd(gnd), .vdd(vdd), .A(_1284_), .Y(_1304_) );
NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_1278_), .B(_1304_), .Y(_1305_) );
OAI21X1 OAI21X1_925 ( .gnd(gnd), .vdd(vdd), .A(_1276_), .B(_1285_), .C(_1305_), .Y(_1306_) );
INVX2 INVX2_54 ( .gnd(gnd), .vdd(vdd), .A(b_reg_25_), .Y(_1307_) );
INVX2 INVX2_55 ( .gnd(gnd), .vdd(vdd), .A(c_reg_25_), .Y(_1308_) );
INVX2 INVX2_56 ( .gnd(gnd), .vdd(vdd), .A(d_reg_25_), .Y(_1309_) );
OAI21X1 OAI21X1_926 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_1307_), .C(_1309_), .Y(_1310_) );
OAI21X1 OAI21X1_927 ( .gnd(gnd), .vdd(vdd), .A(c_reg_25_), .B(_1307_), .C(_1310_), .Y(_1311_) );
NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf4), .B(_1311_), .Y(_1312_) );
NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_1307_), .Y(_1313_) );
NAND3X1 NAND3X1_277 ( .gnd(gnd), .vdd(vdd), .A(_1310_), .B(_1313_), .C(_3451__bF_buf2), .Y(_1314_) );
NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(c_reg_25_), .B(b_reg_25_), .Y(_1315_) );
NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1315_), .B(_1313_), .Y(_1316_) );
XNOR2X1 XNOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1316_), .B(d_reg_25_), .Y(_1317_) );
AOI21X1 AOI21X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1317_), .B(_3405__bF_buf3), .C(_3447__bF_buf3), .Y(_1318_) );
NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(_1314_), .B(_1318_), .Y(_1319_) );
NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1319_), .Y(_1320_) );
AOI21X1 AOI21X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1283_), .B(w_24_), .C(_1281_), .Y(_1321_) );
XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(a_reg_20_), .B(e_reg_25_), .Y(_1322_) );
XNOR2X1 XNOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1322_), .B(w_25_), .Y(_1323_) );
XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_1323_), .B(_1321_), .Y(_1324_) );
XNOR2X1 XNOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1320_), .B(_1324_), .Y(_1325_) );
XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1306_), .Y(_1326_) );
XNOR2X1 XNOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_1326_), .Y(_1327_) );
OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(_1327_), .B(_1302_), .Y(_1328_) );
OAI21X1 OAI21X1_928 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1296_), .C(_1327_), .Y(_1329_) );
OAI21X1 OAI21X1_929 ( .gnd(gnd), .vdd(vdd), .A(_1296_), .B(_1328_), .C(_1329_), .Y(_1330_) );
INVX1 INVX1_706 ( .gnd(gnd), .vdd(vdd), .A(_3667__153_), .Y(_1331_) );
OAI21X1 OAI21X1_930 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1331_), .Y(_1332_) );
AOI22X1 AOI22X1_662 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf10), .B(_1332_), .C(a_reg_25_), .D(_113__bF_buf3), .Y(_1333_) );
OAI21X1 OAI21X1_931 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_1330_), .C(_1333_), .Y(_5__25_) );
INVX1 INVX1_707 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .Y(_1334_) );
INVX1 INVX1_708 ( .gnd(gnd), .vdd(vdd), .A(_1294_), .Y(_1335_) );
OAI21X1 OAI21X1_932 ( .gnd(gnd), .vdd(vdd), .A(_1292_), .B(_1335_), .C(_1327_), .Y(_1336_) );
INVX1 INVX1_709 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .Y(_1337_) );
NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(_1337_), .Y(_1338_) );
NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(_1337_), .Y(_1339_) );
AOI21X1 AOI21X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1302_), .B(_1339_), .C(_1338_), .Y(_1340_) );
OAI21X1 OAI21X1_933 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1334_), .C(_1340_), .Y(_1341_) );
OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(_1325_), .B(_1306_), .Y(_1342_) );
INVX1 INVX1_710 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .Y(_1343_) );
NAND3X1 NAND3X1_278 ( .gnd(gnd), .vdd(vdd), .A(_1312_), .B(_1319_), .C(_1324_), .Y(_1344_) );
OAI21X1 OAI21X1_934 ( .gnd(gnd), .vdd(vdd), .A(_1321_), .B(_1323_), .C(_1344_), .Y(_1345_) );
INVX2 INVX2_57 ( .gnd(gnd), .vdd(vdd), .A(c_reg_26_), .Y(_1346_) );
INVX2 INVX2_58 ( .gnd(gnd), .vdd(vdd), .A(b_reg_26_), .Y(_1347_) );
INVX1 INVX1_711 ( .gnd(gnd), .vdd(vdd), .A(d_reg_26_), .Y(_1348_) );
OAI21X1 OAI21X1_935 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_1347_), .C(_1348_), .Y(_1349_) );
OAI21X1 OAI21X1_936 ( .gnd(gnd), .vdd(vdd), .A(c_reg_26_), .B(b_reg_26_), .C(_1349_), .Y(_1350_) );
XNOR2X1 XNOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(c_reg_26_), .B(b_reg_26_), .Y(_1351_) );
XNOR2X1 XNOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1351_), .B(d_reg_26_), .Y(_1352_) );
OAI21X1 OAI21X1_937 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf1), .B(_40__bF_buf2), .C(_1352_), .Y(_1353_) );
OAI21X1 OAI21X1_938 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf2), .B(_1350_), .C(_1353_), .Y(_1354_) );
OAI21X1 OAI21X1_939 ( .gnd(gnd), .vdd(vdd), .A(c_reg_26_), .B(_1347_), .C(_1349_), .Y(_1355_) );
NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf2), .B(_1355_), .Y(_1356_) );
OAI21X1 OAI21X1_940 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf1), .B(_1354_), .C(_1356_), .Y(_1357_) );
INVX1 INVX1_712 ( .gnd(gnd), .vdd(vdd), .A(a_reg_20_), .Y(_1358_) );
INVX1 INVX1_713 ( .gnd(gnd), .vdd(vdd), .A(e_reg_25_), .Y(_1359_) );
NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(w_25_), .B(_1322_), .Y(_1360_) );
OAI21X1 OAI21X1_941 ( .gnd(gnd), .vdd(vdd), .A(_1358_), .B(_1359_), .C(_1360_), .Y(_1361_) );
INVX1 INVX1_714 ( .gnd(gnd), .vdd(vdd), .A(a_reg_21_), .Y(_1362_) );
INVX1 INVX1_715 ( .gnd(gnd), .vdd(vdd), .A(e_reg_26_), .Y(_1363_) );
NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_1362_), .B(_1363_), .Y(_1364_) );
NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(a_reg_21_), .B(e_reg_26_), .Y(_1365_) );
NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(_1365_), .B(_1364_), .Y(_1366_) );
XNOR2X1 XNOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(w_26_), .Y(_1367_) );
XNOR2X1 XNOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .B(_1361_), .Y(_1368_) );
XNOR2X1 XNOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1357_), .B(_1368_), .Y(_1369_) );
NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1345_), .B(_1369_), .Y(_1370_) );
OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1345_), .Y(_1371_) );
NAND3X1 NAND3X1_279 ( .gnd(gnd), .vdd(vdd), .A(_785_), .B(_1370_), .C(_1371_), .Y(_1372_) );
XNOR2X1 XNOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1369_), .B(_1345_), .Y(_1373_) );
NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_1373_), .Y(_1374_) );
NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(_1372_), .B(_1374_), .Y(_1375_) );
NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1375_), .Y(_1376_) );
NAND3X1 NAND3X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1342_), .B(_1372_), .C(_1374_), .Y(_1377_) );
AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(_1376_), .B(_1377_), .Y(_1378_) );
AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1378_), .Y(_1379_) );
OAI21X1 OAI21X1_942 ( .gnd(gnd), .vdd(vdd), .A(_1378_), .B(_1341_), .C(round_ctr_inc_bF_buf3), .Y(_1380_) );
INVX1 INVX1_716 ( .gnd(gnd), .vdd(vdd), .A(_3667__154_), .Y(_1381_) );
OAI21X1 OAI21X1_943 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1381_), .Y(_1382_) );
AOI22X1 AOI22X1_663 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf9), .B(_1382_), .C(a_reg_26_), .D(_113__bF_buf2), .Y(_1383_) );
OAI21X1 OAI21X1_944 ( .gnd(gnd), .vdd(vdd), .A(_1379_), .B(_1380_), .C(_1383_), .Y(_5__26_) );
INVX1 INVX1_717 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .Y(_1384_) );
AOI21X1 AOI21X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1341_), .B(_1378_), .C(_1384_), .Y(_1385_) );
OAI21X1 OAI21X1_945 ( .gnd(gnd), .vdd(vdd), .A(_786_), .B(_1373_), .C(_1370_), .Y(_1386_) );
INVX1 INVX1_718 ( .gnd(gnd), .vdd(vdd), .A(_1367_), .Y(_1387_) );
NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_1361_), .B(_1387_), .Y(_1388_) );
NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(_1361_), .B(_1387_), .Y(_1389_) );
OAI21X1 OAI21X1_946 ( .gnd(gnd), .vdd(vdd), .A(_1389_), .B(_1357_), .C(_1388_), .Y(_1390_) );
INVX1 INVX1_719 ( .gnd(gnd), .vdd(vdd), .A(c_reg_27_), .Y(_1391_) );
INVX1 INVX1_720 ( .gnd(gnd), .vdd(vdd), .A(b_reg_27_), .Y(_1392_) );
OAI21X1 OAI21X1_947 ( .gnd(gnd), .vdd(vdd), .A(c_reg_27_), .B(b_reg_27_), .C(d_reg_27_), .Y(_1393_) );
OAI21X1 OAI21X1_948 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1392_), .C(_1393_), .Y(_1394_) );
NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(c_reg_27_), .B(b_reg_27_), .Y(_1395_) );
NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(b_reg_27_), .B(d_reg_27_), .Y(_1396_) );
NAND3X1 NAND3X1_281 ( .gnd(gnd), .vdd(vdd), .A(c_reg_27_), .B(b_reg_27_), .C(d_reg_27_), .Y(_1397_) );
AOI22X1 AOI22X1_664 ( .gnd(gnd), .vdd(vdd), .A(_1395_), .B(_1396_), .C(_1397_), .D(_1394_), .Y(_1398_) );
AOI22X1 AOI22X1_665 ( .gnd(gnd), .vdd(vdd), .A(_3451__bF_buf1), .B(_1394_), .C(_1398_), .D(_3474__bF_buf0), .Y(_1399_) );
OAI21X1 OAI21X1_949 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_6_), .B(_3402_), .C(_1399_), .Y(_1400_) );
NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(c_reg_27_), .B(_1392_), .Y(_1401_) );
OAI21X1 OAI21X1_950 ( .gnd(gnd), .vdd(vdd), .A(_1396_), .B(_1401_), .C(_3447__bF_buf0), .Y(_1402_) );
NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_1402_), .B(_1400_), .Y(_1403_) );
AOI21X1 AOI21X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1366_), .B(w_26_), .C(_1364_), .Y(_1404_) );
INVX2 INVX2_59 ( .gnd(gnd), .vdd(vdd), .A(a_reg_22_), .Y(_1405_) );
INVX2 INVX2_60 ( .gnd(gnd), .vdd(vdd), .A(e_reg_27_), .Y(_1406_) );
NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .B(_1406_), .Y(_1407_) );
NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(a_reg_22_), .B(e_reg_27_), .Y(_1408_) );
NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_1408_), .B(_1407_), .Y(_1409_) );
XNOR2X1 XNOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1409_), .B(w_27_), .Y(_1410_) );
XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_1410_), .B(_1404_), .Y(_1411_) );
XNOR2X1 XNOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1403_), .B(_1411_), .Y(_1412_) );
OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(_1412_), .B(_1390_), .Y(_1413_) );
NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1412_), .Y(_1414_) );
NAND3X1 NAND3X1_282 ( .gnd(gnd), .vdd(vdd), .A(_1413_), .B(_1414_), .C(_1386_), .Y(_1415_) );
NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(_1414_), .B(_1413_), .Y(_1416_) );
NAND3X1 NAND3X1_283 ( .gnd(gnd), .vdd(vdd), .A(_1370_), .B(_1416_), .C(_1372_), .Y(_1417_) );
NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_1417_), .B(_1415_), .Y(_1418_) );
INVX1 INVX1_721 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .Y(_1419_) );
AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(_1385_), .B(_1419_), .Y(_1420_) );
OAI21X1 OAI21X1_951 ( .gnd(gnd), .vdd(vdd), .A(_1419_), .B(_1385_), .C(round_ctr_inc_bF_buf2), .Y(_1421_) );
INVX1 INVX1_722 ( .gnd(gnd), .vdd(vdd), .A(_3667__155_), .Y(_1422_) );
NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_3432__bF_buf3), .Y(_1423_) );
AOI22X1 AOI22X1_666 ( .gnd(gnd), .vdd(vdd), .A(_1423_), .B(_3433__bF_buf8), .C(a_reg_27_), .D(_113__bF_buf1), .Y(_1424_) );
OAI21X1 OAI21X1_952 ( .gnd(gnd), .vdd(vdd), .A(_1420_), .B(_1421_), .C(_1424_), .Y(_5__27_) );
NAND3X1 NAND3X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1377_), .B(_1376_), .C(_1418_), .Y(_1425_) );
NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_1336_), .B(_1425_), .Y(_1426_) );
NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1416_), .B(_1386_), .Y(_1427_) );
OAI21X1 OAI21X1_953 ( .gnd(gnd), .vdd(vdd), .A(_1343_), .B(_1375_), .C(_1427_), .Y(_1428_) );
OAI21X1 OAI21X1_954 ( .gnd(gnd), .vdd(vdd), .A(_1386_), .B(_1416_), .C(_1428_), .Y(_1429_) );
OAI21X1 OAI21X1_955 ( .gnd(gnd), .vdd(vdd), .A(_1340_), .B(_1425_), .C(_1429_), .Y(_1430_) );
AOI21X1 AOI21X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1261_), .B(_1426_), .C(_1430_), .Y(_1431_) );
NAND3X1 NAND3X1_285 ( .gnd(gnd), .vdd(vdd), .A(_1400_), .B(_1402_), .C(_1411_), .Y(_1432_) );
OAI21X1 OAI21X1_956 ( .gnd(gnd), .vdd(vdd), .A(_1404_), .B(_1410_), .C(_1432_), .Y(_1433_) );
INVX2 INVX2_61 ( .gnd(gnd), .vdd(vdd), .A(c_reg_28_), .Y(_1434_) );
INVX1 INVX1_723 ( .gnd(gnd), .vdd(vdd), .A(b_reg_28_), .Y(_1435_) );
INVX2 INVX2_62 ( .gnd(gnd), .vdd(vdd), .A(d_reg_28_), .Y(_1436_) );
OAI21X1 OAI21X1_957 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1435_), .C(_1436_), .Y(_1437_) );
OAI21X1 OAI21X1_958 ( .gnd(gnd), .vdd(vdd), .A(c_reg_28_), .B(b_reg_28_), .C(_1437_), .Y(_1438_) );
XNOR2X1 XNOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(c_reg_28_), .B(b_reg_28_), .Y(_1439_) );
XNOR2X1 XNOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1439_), .B(d_reg_28_), .Y(_1440_) );
OAI21X1 OAI21X1_959 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf0), .B(_40__bF_buf1), .C(_1440_), .Y(_1441_) );
OAI21X1 OAI21X1_960 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf1), .B(_1438_), .C(_1441_), .Y(_1442_) );
OAI21X1 OAI21X1_961 ( .gnd(gnd), .vdd(vdd), .A(c_reg_28_), .B(_1435_), .C(_1437_), .Y(_1443_) );
NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf4), .B(_1443_), .Y(_1444_) );
OAI21X1 OAI21X1_962 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf3), .B(_1442_), .C(_1444_), .Y(_1445_) );
NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(w_27_), .B(_1409_), .Y(_1446_) );
OAI21X1 OAI21X1_963 ( .gnd(gnd), .vdd(vdd), .A(_1405_), .B(_1406_), .C(_1446_), .Y(_1447_) );
XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(a_reg_23_), .B(e_reg_28_), .Y(_1448_) );
XNOR2X1 XNOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1448_), .B(w_28_), .Y(_1449_) );
INVX1 INVX1_724 ( .gnd(gnd), .vdd(vdd), .A(_1449_), .Y(_1450_) );
NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1450_), .Y(_1451_) );
INVX1 INVX1_725 ( .gnd(gnd), .vdd(vdd), .A(_1451_), .Y(_1452_) );
NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_1447_), .B(_1450_), .Y(_1453_) );
NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1452_), .Y(_1454_) );
XNOR2X1 XNOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1454_), .B(_1445_), .Y(_1455_) );
OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(_1455_), .B(_1433_), .Y(_1456_) );
NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1433_), .B(_1455_), .Y(_1457_) );
AOI21X1 AOI21X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1456_), .B(_1457_), .C(_3447__bF_buf2), .Y(_1458_) );
NAND3X1 NAND3X1_286 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf1), .B(_1457_), .C(_1456_), .Y(_1459_) );
INVX1 INVX1_726 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .Y(_1460_) );
NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(_1458_), .B(_1460_), .Y(_1461_) );
OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(_1461_), .B(_1413_), .Y(_1462_) );
OAI21X1 OAI21X1_964 ( .gnd(gnd), .vdd(vdd), .A(_1390_), .B(_1412_), .C(_1461_), .Y(_1463_) );
NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .B(_1462_), .Y(_1464_) );
AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(_1431_), .B(_1464_), .Y(_1465_) );
OAI21X1 OAI21X1_965 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1431_), .C(round_ctr_inc_bF_buf1), .Y(_1466_) );
INVX1 INVX1_727 ( .gnd(gnd), .vdd(vdd), .A(_3667__156_), .Y(_1467_) );
NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .B(_3432__bF_buf2), .Y(_1468_) );
AOI22X1 AOI22X1_667 ( .gnd(gnd), .vdd(vdd), .A(_1468_), .B(_3433__bF_buf7), .C(a_reg_28_), .D(_113__bF_buf0), .Y(_1469_) );
OAI21X1 OAI21X1_966 ( .gnd(gnd), .vdd(vdd), .A(_1465_), .B(_1466_), .C(_1469_), .Y(_5__28_) );
AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(_1459_), .B(_1457_), .Y(_1470_) );
OAI21X1 OAI21X1_967 ( .gnd(gnd), .vdd(vdd), .A(_1453_), .B(_1445_), .C(_1451_), .Y(_1471_) );
INVX2 INVX2_63 ( .gnd(gnd), .vdd(vdd), .A(b_reg_29_), .Y(_1472_) );
INVX1 INVX1_728 ( .gnd(gnd), .vdd(vdd), .A(c_reg_29_), .Y(_1473_) );
INVX2 INVX2_64 ( .gnd(gnd), .vdd(vdd), .A(d_reg_29_), .Y(_1474_) );
OAI21X1 OAI21X1_968 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(_1472_), .C(_1474_), .Y(_1475_) );
OAI21X1 OAI21X1_969 ( .gnd(gnd), .vdd(vdd), .A(c_reg_29_), .B(_1472_), .C(_1475_), .Y(_1476_) );
NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf0), .B(_1476_), .Y(_1477_) );
OAI21X1 OAI21X1_970 ( .gnd(gnd), .vdd(vdd), .A(c_reg_29_), .B(b_reg_29_), .C(_1475_), .Y(_1478_) );
XNOR2X1 XNOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(c_reg_29_), .B(b_reg_29_), .Y(_1479_) );
XNOR2X1 XNOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1479_), .B(_1474_), .Y(_1480_) );
OAI22X1 OAI22X1_60 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf0), .B(_1478_), .C(_3406__bF_buf2), .D(_1480_), .Y(_1481_) );
OAI21X1 OAI21X1_971 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf4), .B(_1481_), .C(_1477_), .Y(_1482_) );
INVX1 INVX1_729 ( .gnd(gnd), .vdd(vdd), .A(a_reg_23_), .Y(_1483_) );
INVX2 INVX2_65 ( .gnd(gnd), .vdd(vdd), .A(e_reg_28_), .Y(_1484_) );
NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(w_28_), .B(_1448_), .Y(_1485_) );
OAI21X1 OAI21X1_972 ( .gnd(gnd), .vdd(vdd), .A(_1483_), .B(_1484_), .C(_1485_), .Y(_1486_) );
INVX1 INVX1_730 ( .gnd(gnd), .vdd(vdd), .A(w_29_), .Y(_1487_) );
INVX2 INVX2_66 ( .gnd(gnd), .vdd(vdd), .A(e_reg_29_), .Y(_1488_) );
NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_1247_), .B(_1488_), .Y(_1489_) );
NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(a_reg_24_), .B(e_reg_29_), .Y(_1490_) );
NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_1490_), .B(_1489_), .Y(_1491_) );
XNOR2X1 XNOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1491_), .B(_1487_), .Y(_1492_) );
XNOR2X1 XNOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1492_), .B(_1486_), .Y(_1493_) );
OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(_1493_), .B(_1482_), .Y(_1494_) );
NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(_1482_), .B(_1493_), .Y(_1495_) );
NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_1495_), .B(_1494_), .Y(_1496_) );
XNOR2X1 XNOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1496_), .B(_1471_), .Y(_1497_) );
XNOR2X1 XNOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1497_), .B(_40__bF_buf0), .Y(_1498_) );
XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_1470_), .B(_1498_), .Y(_1499_) );
OAI21X1 OAI21X1_973 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1431_), .C(_1463_), .Y(_1500_) );
XNOR2X1 XNOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1500_), .B(_1499_), .Y(_1501_) );
INVX1 INVX1_731 ( .gnd(gnd), .vdd(vdd), .A(_3667__157_), .Y(_1502_) );
OAI21X1 OAI21X1_974 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1502_), .Y(_1503_) );
AOI22X1 AOI22X1_668 ( .gnd(gnd), .vdd(vdd), .A(_3433__bF_buf6), .B(_1503_), .C(a_reg_29_), .D(_113__bF_buf4), .Y(_1504_) );
OAI21X1 OAI21X1_975 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_1501_), .C(_1504_), .Y(_5__29_) );
NAND3X1 NAND3X1_287 ( .gnd(gnd), .vdd(vdd), .A(_1184_), .B(_1133_), .C(_1241_), .Y(_1505_) );
NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_1018_), .B(_1505_), .Y(_1506_) );
OAI21X1 OAI21X1_976 ( .gnd(gnd), .vdd(vdd), .A(_782_), .B(_776_), .C(_1506_), .Y(_1507_) );
NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_1326_), .B(_1303_), .Y(_1508_) );
OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(_1303_), .B(_1326_), .Y(_1509_) );
AOI22X1 AOI22X1_669 ( .gnd(gnd), .vdd(vdd), .A(_1508_), .B(_1509_), .C(_1294_), .D(_1293_), .Y(_1510_) );
NAND3X1 NAND3X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1418_), .B(_1378_), .C(_1510_), .Y(_1511_) );
AOI21X1 AOI21X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1507_), .B(_1260_), .C(_1511_), .Y(_1512_) );
INVX1 INVX1_732 ( .gnd(gnd), .vdd(vdd), .A(_1499_), .Y(_1513_) );
NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_1513_), .B(_1464_), .Y(_1514_) );
OAI21X1 OAI21X1_977 ( .gnd(gnd), .vdd(vdd), .A(_1430_), .B(_1512_), .C(_1514_), .Y(_1515_) );
INVX1 INVX1_733 ( .gnd(gnd), .vdd(vdd), .A(_1463_), .Y(_1516_) );
NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(_1498_), .B(_1470_), .Y(_1517_) );
AOI21X1 AOI21X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1516_), .B(_1499_), .C(_1517_), .Y(_1518_) );
NAND3X1 NAND3X1_289 ( .gnd(gnd), .vdd(vdd), .A(_1494_), .B(_1495_), .C(_1471_), .Y(_1519_) );
NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_40__bF_buf3), .B(_1497_), .Y(_1520_) );
NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(_1519_), .B(_1520_), .Y(_1521_) );
NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_1486_), .B(_1492_), .Y(_1522_) );
OAI21X1 OAI21X1_978 ( .gnd(gnd), .vdd(vdd), .A(_1482_), .B(_1493_), .C(_1522_), .Y(_1523_) );
INVX2 INVX2_67 ( .gnd(gnd), .vdd(vdd), .A(c_reg_30_), .Y(_1524_) );
INVX1 INVX1_734 ( .gnd(gnd), .vdd(vdd), .A(b_reg_30_), .Y(_1525_) );
INVX1 INVX1_735 ( .gnd(gnd), .vdd(vdd), .A(d_reg_30_), .Y(_1526_) );
OAI21X1 OAI21X1_979 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1525_), .C(_1526_), .Y(_1527_) );
OAI21X1 OAI21X1_980 ( .gnd(gnd), .vdd(vdd), .A(c_reg_30_), .B(b_reg_30_), .C(_1527_), .Y(_1528_) );
XNOR2X1 XNOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(c_reg_30_), .B(b_reg_30_), .Y(_1529_) );
XNOR2X1 XNOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1529_), .B(d_reg_30_), .Y(_1530_) );
OAI21X1 OAI21X1_981 ( .gnd(gnd), .vdd(vdd), .A(_3437__bF_buf3), .B(_40__bF_buf2), .C(_1530_), .Y(_1531_) );
OAI21X1 OAI21X1_982 ( .gnd(gnd), .vdd(vdd), .A(_3405__bF_buf5), .B(_1528_), .C(_1531_), .Y(_1532_) );
OAI21X1 OAI21X1_983 ( .gnd(gnd), .vdd(vdd), .A(c_reg_30_), .B(_1525_), .C(_1527_), .Y(_1533_) );
NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf3), .B(_1533_), .Y(_1534_) );
OAI21X1 OAI21X1_984 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf2), .B(_1532_), .C(_1534_), .Y(_1535_) );
INVX1 INVX1_736 ( .gnd(gnd), .vdd(vdd), .A(_1489_), .Y(_1536_) );
OAI21X1 OAI21X1_985 ( .gnd(gnd), .vdd(vdd), .A(_1487_), .B(_1490_), .C(_1536_), .Y(_1537_) );
INVX1 INVX1_737 ( .gnd(gnd), .vdd(vdd), .A(a_reg_25_), .Y(_1538_) );
INVX1 INVX1_738 ( .gnd(gnd), .vdd(vdd), .A(e_reg_30_), .Y(_1539_) );
NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1539_), .Y(_1540_) );
NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(a_reg_25_), .B(e_reg_30_), .Y(_1541_) );
NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(_1541_), .B(_1540_), .Y(_1542_) );
NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(w_30_), .B(_1542_), .Y(_1543_) );
OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(_1542_), .B(w_30_), .Y(_1544_) );
AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(_1544_), .B(_1543_), .Y(_1545_) );
XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_1545_), .B(_1537_), .Y(_1546_) );
XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(_1546_), .Y(_1547_) );
XNOR2X1 XNOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1547_), .B(_1523_), .Y(_1548_) );
XNOR2X1 XNOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1548_), .B(_3405__bF_buf4), .Y(_1549_) );
OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(_1549_), .B(_1521_), .Y(_1550_) );
NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_1521_), .B(_1549_), .Y(_1551_) );
AOI22X1 AOI22X1_670 ( .gnd(gnd), .vdd(vdd), .A(_1550_), .B(_1551_), .C(_1518_), .D(_1515_), .Y(_1552_) );
OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(_1464_), .B(_1513_), .Y(_1553_) );
OAI21X1 OAI21X1_986 ( .gnd(gnd), .vdd(vdd), .A(_1553_), .B(_1431_), .C(_1518_), .Y(_1554_) );
NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(_1551_), .B(_1550_), .Y(_1555_) );
OAI21X1 OAI21X1_987 ( .gnd(gnd), .vdd(vdd), .A(_1555_), .B(_1554_), .C(round_ctr_inc_bF_buf0), .Y(_1556_) );
OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(_3432__bF_buf1), .B(_3667__158_), .Y(_1557_) );
AOI22X1 AOI22X1_671 ( .gnd(gnd), .vdd(vdd), .A(_113__bF_buf3), .B(a_reg_30_), .C(_3433__bF_buf5), .D(_1557_), .Y(_1558_) );
OAI21X1 OAI21X1_988 ( .gnd(gnd), .vdd(vdd), .A(_1552_), .B(_1556_), .C(_1558_), .Y(_5__30_) );
AOI21X1 AOI21X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1519_), .B(_1520_), .C(_1549_), .Y(_1559_) );
INVX1 INVX1_739 ( .gnd(gnd), .vdd(vdd), .A(_1523_), .Y(_1560_) );
OAI21X1 OAI21X1_989 ( .gnd(gnd), .vdd(vdd), .A(_3392_), .B(_3437__bF_buf2), .C(_1548_), .Y(_1561_) );
OAI21X1 OAI21X1_990 ( .gnd(gnd), .vdd(vdd), .A(_1560_), .B(_1547_), .C(_1561_), .Y(_1562_) );
NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_1537_), .B(_1545_), .Y(_1563_) );
INVX1 INVX1_740 ( .gnd(gnd), .vdd(vdd), .A(_1546_), .Y(_1564_) );
OAI21X1 OAI21X1_991 ( .gnd(gnd), .vdd(vdd), .A(_1535_), .B(_1564_), .C(_1563_), .Y(_1565_) );
INVX1 INVX1_741 ( .gnd(gnd), .vdd(vdd), .A(c_reg_31_), .Y(_1566_) );
INVX1 INVX1_742 ( .gnd(gnd), .vdd(vdd), .A(b_reg_31_), .Y(_1567_) );
OAI21X1 OAI21X1_992 ( .gnd(gnd), .vdd(vdd), .A(c_reg_31_), .B(b_reg_31_), .C(d_reg_31_), .Y(_1568_) );
OAI21X1 OAI21X1_993 ( .gnd(gnd), .vdd(vdd), .A(_1566_), .B(_1567_), .C(_1568_), .Y(_1569_) );
NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(_1569_), .B(_3451__bF_buf0), .Y(_1570_) );
NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_1566_), .B(_1567_), .Y(_1571_) );
NAND3X1 NAND3X1_290 ( .gnd(gnd), .vdd(vdd), .A(c_reg_31_), .B(b_reg_31_), .C(d_reg_31_), .Y(_1572_) );
NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(_1572_), .B(_1569_), .Y(_1573_) );
OAI21X1 OAI21X1_994 ( .gnd(gnd), .vdd(vdd), .A(d_reg_31_), .B(_1571_), .C(_1573_), .Y(_1574_) );
OAI21X1 OAI21X1_995 ( .gnd(gnd), .vdd(vdd), .A(_3406__bF_buf1), .B(_1574_), .C(_1570_), .Y(_1575_) );
NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(b_reg_31_), .B(d_reg_31_), .Y(_1576_) );
NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(c_reg_31_), .B(_1567_), .Y(_1577_) );
OAI21X1 OAI21X1_996 ( .gnd(gnd), .vdd(vdd), .A(_1576_), .B(_1577_), .C(_3447__bF_buf1), .Y(_1578_) );
OAI21X1 OAI21X1_997 ( .gnd(gnd), .vdd(vdd), .A(_3447__bF_buf0), .B(_1575_), .C(_1578_), .Y(_1579_) );
OAI21X1 OAI21X1_998 ( .gnd(gnd), .vdd(vdd), .A(_1538_), .B(_1539_), .C(_1543_), .Y(_1580_) );
XNOR2X1 XNOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(a_reg_26_), .B(w_31_), .Y(_1581_) );
XNOR2X1 XNOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1581_), .B(e_reg_31_), .Y(_1582_) );
XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_1580_), .B(_1582_), .Y(_1583_) );
XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_1583_), .B(_1579_), .Y(_1584_) );
XNOR2X1 XNOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(_1565_), .B(_1584_), .Y(_1585_) );
XNOR2X1 XNOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(_1585_), .B(_3392_), .Y(_1586_) );
XNOR2X1 XNOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(_1562_), .B(_1586_), .Y(_1587_) );
INVX1 INVX1_743 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .Y(_1588_) );
NOR3X1 NOR3X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1559_), .B(_1588_), .C(_1552_), .Y(_1589_) );
AOI21X1 AOI21X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1554_), .B(_1555_), .C(_1559_), .Y(_1590_) );
OAI21X1 OAI21X1_999 ( .gnd(gnd), .vdd(vdd), .A(_1587_), .B(_1590_), .C(round_ctr_inc_bF_buf11), .Y(_1591_) );
INVX1 INVX1_744 ( .gnd(gnd), .vdd(vdd), .A(_3667__159_), .Y(_1592_) );
NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_1592_), .B(_3432__bF_buf0), .Y(_1593_) );
AOI22X1 AOI22X1_672 ( .gnd(gnd), .vdd(vdd), .A(_1593_), .B(_3433__bF_buf4), .C(a_reg_31_), .D(_113__bF_buf2), .Y(_1594_) );
OAI21X1 OAI21X1_1000 ( .gnd(gnd), .vdd(vdd), .A(_1589_), .B(_1591_), .C(_1594_), .Y(_5__31_) );
INVX1 INVX1_745 ( .gnd(gnd), .vdd(vdd), .A(_3667__96_), .Y(_1595_) );
OAI21X1 OAI21X1_1001 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1595_), .Y(_1596_) );
AOI22X1 AOI22X1_673 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(a_reg_0_), .C(_1596_), .D(_3433__bF_buf3), .Y(_1597_) );
OAI21X1 OAI21X1_1002 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_3387__bF_buf0), .C(_1597_), .Y(_6__0_) );
INVX1 INVX1_746 ( .gnd(gnd), .vdd(vdd), .A(_3667__97_), .Y(_1598_) );
NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .B(_3432__bF_buf11), .Y(_1599_) );
AOI22X1 AOI22X1_674 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(a_reg_1_), .C(_3433__bF_buf2), .D(_1599_), .Y(_1600_) );
OAI21X1 OAI21X1_1003 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_3387__bF_buf10), .C(_1600_), .Y(_6__1_) );
INVX1 INVX1_747 ( .gnd(gnd), .vdd(vdd), .A(b_reg_2_), .Y(_1601_) );
INVX1 INVX1_748 ( .gnd(gnd), .vdd(vdd), .A(_3667__98_), .Y(_1602_) );
NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_3432__bF_buf10), .Y(_1603_) );
AOI22X1 AOI22X1_675 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(a_reg_2_), .C(_3433__bF_buf1), .D(_1603_), .Y(_1604_) );
OAI21X1 OAI21X1_1004 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .B(_3387__bF_buf9), .C(_1604_), .Y(_6__2_) );
INVX1 INVX1_749 ( .gnd(gnd), .vdd(vdd), .A(_3667__99_), .Y(_1605_) );
OAI21X1 OAI21X1_1005 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1605_), .Y(_1606_) );
AOI22X1 AOI22X1_676 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(a_reg_3_), .C(_1606_), .D(_3433__bF_buf0), .Y(_1607_) );
OAI21X1 OAI21X1_1006 ( .gnd(gnd), .vdd(vdd), .A(_3575_), .B(_3387__bF_buf8), .C(_1607_), .Y(_6__3_) );
INVX1 INVX1_750 ( .gnd(gnd), .vdd(vdd), .A(_3667__100_), .Y(_1608_) );
NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_3432__bF_buf9), .Y(_1609_) );
AOI22X1 AOI22X1_677 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(a_reg_4_), .C(_3433__bF_buf11), .D(_1609_), .Y(_1610_) );
OAI21X1 OAI21X1_1007 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_3387__bF_buf7), .C(_1610_), .Y(_6__4_) );
INVX1 INVX1_751 ( .gnd(gnd), .vdd(vdd), .A(_3667__101_), .Y(_1611_) );
NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_3432__bF_buf8), .Y(_1612_) );
AOI22X1 AOI22X1_678 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(a_reg_5_), .C(_3433__bF_buf10), .D(_1612_), .Y(_1613_) );
OAI21X1 OAI21X1_1008 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_3387__bF_buf6), .C(_1613_), .Y(_6__5_) );
INVX1 INVX1_752 ( .gnd(gnd), .vdd(vdd), .A(b_reg_6_), .Y(_1614_) );
INVX2 INVX2_68 ( .gnd(gnd), .vdd(vdd), .A(_3667__102_), .Y(_1615_) );
NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_3432__bF_buf7), .Y(_1616_) );
AOI22X1 AOI22X1_679 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(a_reg_6_), .C(_3433__bF_buf9), .D(_1616_), .Y(_1617_) );
OAI21X1 OAI21X1_1009 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .B(_3387__bF_buf5), .C(_1617_), .Y(_6__6_) );
OAI21X1 OAI21X1_1010 ( .gnd(gnd), .vdd(vdd), .A(_3667__103_), .B(_3432__bF_buf6), .C(_3433__bF_buf8), .Y(_1618_) );
AOI22X1 AOI22X1_680 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(a_reg_7_), .C(b_reg_7_), .D(_113__bF_buf1), .Y(_1619_) );
NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_1618_), .B(_1619_), .Y(_6__7_) );
INVX1 INVX1_753 ( .gnd(gnd), .vdd(vdd), .A(b_reg_8_), .Y(_1620_) );
INVX1 INVX1_754 ( .gnd(gnd), .vdd(vdd), .A(_3667__104_), .Y(_1621_) );
OAI21X1 OAI21X1_1011 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1621_), .Y(_1622_) );
AOI22X1 AOI22X1_681 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(a_reg_8_), .C(_1622_), .D(_3433__bF_buf7), .Y(_1623_) );
OAI21X1 OAI21X1_1012 ( .gnd(gnd), .vdd(vdd), .A(_1620_), .B(_3387__bF_buf4), .C(_1623_), .Y(_6__8_) );
INVX1 INVX1_755 ( .gnd(gnd), .vdd(vdd), .A(_3667__105_), .Y(_1624_) );
OAI21X1 OAI21X1_1013 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1624_), .Y(_1625_) );
AOI22X1 AOI22X1_682 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(a_reg_9_), .C(_1625_), .D(_3433__bF_buf6), .Y(_1626_) );
OAI21X1 OAI21X1_1014 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_3387__bF_buf3), .C(_1626_), .Y(_6__9_) );
INVX1 INVX1_756 ( .gnd(gnd), .vdd(vdd), .A(b_reg_10_), .Y(_1627_) );
INVX1 INVX1_757 ( .gnd(gnd), .vdd(vdd), .A(_3667__106_), .Y(_1628_) );
NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(_1628_), .B(_3432__bF_buf5), .Y(_1629_) );
AOI22X1 AOI22X1_683 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(a_reg_10_), .C(_3433__bF_buf5), .D(_1629_), .Y(_1630_) );
OAI21X1 OAI21X1_1015 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(_3387__bF_buf2), .C(_1630_), .Y(_6__10_) );
INVX1 INVX1_758 ( .gnd(gnd), .vdd(vdd), .A(b_reg_11_), .Y(_1631_) );
INVX1 INVX1_759 ( .gnd(gnd), .vdd(vdd), .A(_3667__107_), .Y(_1632_) );
OAI21X1 OAI21X1_1016 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1632_), .Y(_1633_) );
AOI22X1 AOI22X1_684 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(a_reg_11_), .C(_1633_), .D(_3433__bF_buf4), .Y(_1634_) );
OAI21X1 OAI21X1_1017 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_3387__bF_buf1), .C(_1634_), .Y(_6__11_) );
INVX1 INVX1_760 ( .gnd(gnd), .vdd(vdd), .A(b_reg_12_), .Y(_1635_) );
INVX1 INVX1_761 ( .gnd(gnd), .vdd(vdd), .A(_3667__108_), .Y(_1636_) );
NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_3432__bF_buf4), .Y(_1637_) );
AOI22X1 AOI22X1_685 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(a_reg_12_), .C(_3433__bF_buf3), .D(_1637_), .Y(_1638_) );
OAI21X1 OAI21X1_1018 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_3387__bF_buf0), .C(_1638_), .Y(_6__12_) );
INVX1 INVX1_762 ( .gnd(gnd), .vdd(vdd), .A(b_reg_13_), .Y(_1639_) );
INVX1 INVX1_763 ( .gnd(gnd), .vdd(vdd), .A(_3667__109_), .Y(_1640_) );
OAI21X1 OAI21X1_1019 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1640_), .Y(_1641_) );
AOI22X1 AOI22X1_686 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(a_reg_13_), .C(_1641_), .D(_3433__bF_buf2), .Y(_1642_) );
OAI21X1 OAI21X1_1020 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_3387__bF_buf10), .C(_1642_), .Y(_6__13_) );
INVX1 INVX1_764 ( .gnd(gnd), .vdd(vdd), .A(b_reg_14_), .Y(_1643_) );
INVX2 INVX2_69 ( .gnd(gnd), .vdd(vdd), .A(_3667__110_), .Y(_1644_) );
NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_1644_), .B(_3432__bF_buf3), .Y(_1645_) );
AOI22X1 AOI22X1_687 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(a_reg_14_), .C(_3433__bF_buf1), .D(_1645_), .Y(_1646_) );
OAI21X1 OAI21X1_1021 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_3387__bF_buf9), .C(_1646_), .Y(_6__14_) );
INVX1 INVX1_765 ( .gnd(gnd), .vdd(vdd), .A(_3667__111_), .Y(_1647_) );
OAI21X1 OAI21X1_1022 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1647_), .Y(_1648_) );
AOI22X1 AOI22X1_688 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(a_reg_15_), .C(_1648_), .D(_3433__bF_buf0), .Y(_1649_) );
OAI21X1 OAI21X1_1023 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_3387__bF_buf8), .C(_1649_), .Y(_6__15_) );
INVX1 INVX1_766 ( .gnd(gnd), .vdd(vdd), .A(_3667__112_), .Y(_1650_) );
OAI21X1 OAI21X1_1024 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1650_), .Y(_1651_) );
AOI22X1 AOI22X1_689 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(a_reg_16_), .C(_1651_), .D(_3433__bF_buf11), .Y(_1652_) );
OAI21X1 OAI21X1_1025 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_3387__bF_buf7), .C(_1652_), .Y(_6__16_) );
INVX1 INVX1_767 ( .gnd(gnd), .vdd(vdd), .A(_3667__113_), .Y(_1653_) );
NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_3432__bF_buf2), .Y(_1654_) );
AOI22X1 AOI22X1_690 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(a_reg_17_), .C(_3433__bF_buf10), .D(_1654_), .Y(_1655_) );
OAI21X1 OAI21X1_1026 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_3387__bF_buf6), .C(_1655_), .Y(_6__17_) );
INVX1 INVX1_768 ( .gnd(gnd), .vdd(vdd), .A(_3667__114_), .Y(_1656_) );
OAI21X1 OAI21X1_1027 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1656_), .Y(_1657_) );
AOI22X1 AOI22X1_691 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(a_reg_18_), .C(_1657_), .D(_3433__bF_buf9), .Y(_1658_) );
OAI21X1 OAI21X1_1028 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_3387__bF_buf5), .C(_1658_), .Y(_6__18_) );
INVX1 INVX1_769 ( .gnd(gnd), .vdd(vdd), .A(_3667__115_), .Y(_1659_) );
OAI21X1 OAI21X1_1029 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1659_), .Y(_1660_) );
AOI22X1 AOI22X1_692 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(a_reg_19_), .C(_1660_), .D(_3433__bF_buf8), .Y(_1661_) );
OAI21X1 OAI21X1_1030 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_3387__bF_buf4), .C(_1661_), .Y(_6__19_) );
INVX1 INVX1_770 ( .gnd(gnd), .vdd(vdd), .A(_3667__116_), .Y(_1662_) );
NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(_1662_), .B(_3432__bF_buf1), .Y(_1663_) );
AOI22X1 AOI22X1_693 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(a_reg_20_), .C(_3433__bF_buf7), .D(_1663_), .Y(_1664_) );
OAI21X1 OAI21X1_1031 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_3387__bF_buf3), .C(_1664_), .Y(_6__20_) );
INVX2 INVX2_70 ( .gnd(gnd), .vdd(vdd), .A(_3667__117_), .Y(_1665_) );
NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_3432__bF_buf0), .Y(_1666_) );
AOI22X1 AOI22X1_694 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(a_reg_21_), .C(_3433__bF_buf6), .D(_1666_), .Y(_1667_) );
OAI21X1 OAI21X1_1032 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_3387__bF_buf2), .C(_1667_), .Y(_6__21_) );
INVX1 INVX1_771 ( .gnd(gnd), .vdd(vdd), .A(_3667__118_), .Y(_1668_) );
OAI21X1 OAI21X1_1033 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1668_), .Y(_1669_) );
AOI22X1 AOI22X1_695 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(a_reg_22_), .C(_1669_), .D(_3433__bF_buf5), .Y(_1670_) );
OAI21X1 OAI21X1_1034 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_3387__bF_buf1), .C(_1670_), .Y(_6__22_) );
INVX1 INVX1_772 ( .gnd(gnd), .vdd(vdd), .A(_3667__119_), .Y(_1671_) );
OAI21X1 OAI21X1_1035 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1671_), .Y(_1672_) );
AOI22X1 AOI22X1_696 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(a_reg_23_), .C(_1672_), .D(_3433__bF_buf4), .Y(_1673_) );
OAI21X1 OAI21X1_1036 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(_3387__bF_buf0), .C(_1673_), .Y(_6__23_) );
INVX1 INVX1_773 ( .gnd(gnd), .vdd(vdd), .A(_3667__120_), .Y(_1674_) );
OAI21X1 OAI21X1_1037 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1674_), .Y(_1675_) );
AOI22X1 AOI22X1_697 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(a_reg_24_), .C(_1675_), .D(_3433__bF_buf3), .Y(_1676_) );
OAI21X1 OAI21X1_1038 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_3387__bF_buf10), .C(_1676_), .Y(_6__24_) );
INVX1 INVX1_774 ( .gnd(gnd), .vdd(vdd), .A(_3667__121_), .Y(_1677_) );
OAI21X1 OAI21X1_1039 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1677_), .Y(_1678_) );
AOI22X1 AOI22X1_698 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(a_reg_25_), .C(_1678_), .D(_3433__bF_buf2), .Y(_1679_) );
OAI21X1 OAI21X1_1040 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_3387__bF_buf9), .C(_1679_), .Y(_6__25_) );
INVX1 INVX1_775 ( .gnd(gnd), .vdd(vdd), .A(_3667__122_), .Y(_1680_) );
OAI21X1 OAI21X1_1041 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1680_), .Y(_1681_) );
AOI22X1 AOI22X1_699 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(a_reg_26_), .C(_1681_), .D(_3433__bF_buf1), .Y(_1682_) );
OAI21X1 OAI21X1_1042 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(_3387__bF_buf8), .C(_1682_), .Y(_6__26_) );
OAI21X1 OAI21X1_1043 ( .gnd(gnd), .vdd(vdd), .A(_3667__123_), .B(_3432__bF_buf11), .C(_3433__bF_buf0), .Y(_1683_) );
AOI22X1 AOI22X1_700 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(a_reg_27_), .C(b_reg_27_), .D(_113__bF_buf0), .Y(_1684_) );
NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(_1683_), .B(_1684_), .Y(_6__27_) );
INVX1 INVX1_776 ( .gnd(gnd), .vdd(vdd), .A(_3667__124_), .Y(_1685_) );
NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_3432__bF_buf10), .Y(_1686_) );
AOI22X1 AOI22X1_701 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(a_reg_28_), .C(_3433__bF_buf11), .D(_1686_), .Y(_1687_) );
OAI21X1 OAI21X1_1044 ( .gnd(gnd), .vdd(vdd), .A(_1435_), .B(_3387__bF_buf7), .C(_1687_), .Y(_6__28_) );
INVX1 INVX1_777 ( .gnd(gnd), .vdd(vdd), .A(_3667__125_), .Y(_1688_) );
OAI21X1 OAI21X1_1045 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1688_), .Y(_1689_) );
AOI22X1 AOI22X1_702 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(a_reg_29_), .C(_1689_), .D(_3433__bF_buf10), .Y(_1690_) );
OAI21X1 OAI21X1_1046 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .B(_3387__bF_buf6), .C(_1690_), .Y(_6__29_) );
OAI21X1 OAI21X1_1047 ( .gnd(gnd), .vdd(vdd), .A(_3667__126_), .B(_3432__bF_buf9), .C(_3433__bF_buf9), .Y(_1691_) );
AOI22X1 AOI22X1_703 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(a_reg_30_), .C(b_reg_30_), .D(_113__bF_buf4), .Y(_1692_) );
NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_1691_), .B(_1692_), .Y(_6__30_) );
OAI21X1 OAI21X1_1048 ( .gnd(gnd), .vdd(vdd), .A(_3667__127_), .B(_3432__bF_buf8), .C(_3433__bF_buf8), .Y(_1693_) );
AOI22X1 AOI22X1_704 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(a_reg_31_), .C(b_reg_31_), .D(_113__bF_buf3), .Y(_1694_) );
NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(_1693_), .B(_1694_), .Y(_6__31_) );
INVX1 INVX1_778 ( .gnd(gnd), .vdd(vdd), .A(_3667__64_), .Y(_1695_) );
NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_3432__bF_buf7), .Y(_1696_) );
AOI22X1 AOI22X1_705 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(b_reg_2_), .C(_3433__bF_buf7), .D(_1696_), .Y(_1697_) );
OAI21X1 OAI21X1_1049 ( .gnd(gnd), .vdd(vdd), .A(_3413_), .B(_3387__bF_buf5), .C(_1697_), .Y(_7__0_) );
INVX1 INVX1_779 ( .gnd(gnd), .vdd(vdd), .A(_3667__65_), .Y(_1698_) );
OAI21X1 OAI21X1_1050 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1698_), .Y(_1699_) );
AOI22X1 AOI22X1_706 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(b_reg_3_), .C(_1699_), .D(_3433__bF_buf6), .Y(_1700_) );
OAI21X1 OAI21X1_1051 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_3387__bF_buf4), .C(_1700_), .Y(_7__1_) );
INVX1 INVX1_780 ( .gnd(gnd), .vdd(vdd), .A(c_reg_2_), .Y(_1701_) );
INVX1 INVX1_781 ( .gnd(gnd), .vdd(vdd), .A(_3667__66_), .Y(_1702_) );
OAI21X1 OAI21X1_1052 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1702_), .Y(_1703_) );
AOI22X1 AOI22X1_707 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(b_reg_4_), .C(_1703_), .D(_3433__bF_buf5), .Y(_1704_) );
OAI21X1 OAI21X1_1053 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(_3387__bF_buf3), .C(_1704_), .Y(_7__2_) );
INVX1 INVX1_782 ( .gnd(gnd), .vdd(vdd), .A(_3667__67_), .Y(_1705_) );
OAI21X1 OAI21X1_1054 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1705_), .Y(_1706_) );
AOI22X1 AOI22X1_708 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(b_reg_5_), .C(_1706_), .D(_3433__bF_buf4), .Y(_1707_) );
OAI21X1 OAI21X1_1055 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_3387__bF_buf2), .C(_1707_), .Y(_7__3_) );
INVX1 INVX1_783 ( .gnd(gnd), .vdd(vdd), .A(_3667__68_), .Y(_1708_) );
OAI21X1 OAI21X1_1056 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1708_), .Y(_1709_) );
AOI22X1 AOI22X1_709 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(b_reg_6_), .C(_1709_), .D(_3433__bF_buf3), .Y(_1710_) );
OAI21X1 OAI21X1_1057 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_3387__bF_buf1), .C(_1710_), .Y(_7__4_) );
INVX1 INVX1_784 ( .gnd(gnd), .vdd(vdd), .A(_3667__69_), .Y(_1711_) );
OAI21X1 OAI21X1_1058 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1711_), .Y(_1712_) );
AOI22X1 AOI22X1_710 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(b_reg_7_), .C(_1712_), .D(_3433__bF_buf2), .Y(_1713_) );
OAI21X1 OAI21X1_1059 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_3387__bF_buf0), .C(_1713_), .Y(_7__5_) );
INVX1 INVX1_785 ( .gnd(gnd), .vdd(vdd), .A(c_reg_6_), .Y(_1714_) );
INVX1 INVX1_786 ( .gnd(gnd), .vdd(vdd), .A(_3667__70_), .Y(_1715_) );
OAI21X1 OAI21X1_1060 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1715_), .Y(_1716_) );
AOI22X1 AOI22X1_711 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(b_reg_8_), .C(_1716_), .D(_3433__bF_buf1), .Y(_1717_) );
OAI21X1 OAI21X1_1061 ( .gnd(gnd), .vdd(vdd), .A(_1714_), .B(_3387__bF_buf10), .C(_1717_), .Y(_7__6_) );
INVX1 INVX1_787 ( .gnd(gnd), .vdd(vdd), .A(_3667__71_), .Y(_1718_) );
OAI21X1 OAI21X1_1062 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1718_), .Y(_1719_) );
AOI22X1 AOI22X1_712 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(b_reg_9_), .C(_1719_), .D(_3433__bF_buf0), .Y(_1720_) );
OAI21X1 OAI21X1_1063 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_3387__bF_buf9), .C(_1720_), .Y(_7__7_) );
INVX1 INVX1_788 ( .gnd(gnd), .vdd(vdd), .A(_3667__72_), .Y(_1721_) );
NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(_3432__bF_buf6), .Y(_1722_) );
AOI22X1 AOI22X1_713 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(b_reg_10_), .C(_3433__bF_buf11), .D(_1722_), .Y(_1723_) );
OAI21X1 OAI21X1_1064 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_3387__bF_buf8), .C(_1723_), .Y(_7__8_) );
INVX2 INVX2_71 ( .gnd(gnd), .vdd(vdd), .A(_3667__73_), .Y(_1724_) );
NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_3432__bF_buf5), .Y(_1725_) );
AOI22X1 AOI22X1_714 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(b_reg_11_), .C(_3433__bF_buf10), .D(_1725_), .Y(_1726_) );
OAI21X1 OAI21X1_1065 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_3387__bF_buf7), .C(_1726_), .Y(_7__9_) );
INVX1 INVX1_789 ( .gnd(gnd), .vdd(vdd), .A(_3667__74_), .Y(_1727_) );
OAI21X1 OAI21X1_1066 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1727_), .Y(_1728_) );
AOI22X1 AOI22X1_715 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(b_reg_12_), .C(_1728_), .D(_3433__bF_buf9), .Y(_1729_) );
OAI21X1 OAI21X1_1067 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_3387__bF_buf6), .C(_1729_), .Y(_7__10_) );
INVX1 INVX1_790 ( .gnd(gnd), .vdd(vdd), .A(_3667__75_), .Y(_1730_) );
OAI21X1 OAI21X1_1068 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1730_), .Y(_1731_) );
AOI22X1 AOI22X1_716 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(b_reg_13_), .C(_1731_), .D(_3433__bF_buf8), .Y(_1732_) );
OAI21X1 OAI21X1_1069 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_3387__bF_buf5), .C(_1732_), .Y(_7__11_) );
INVX1 INVX1_791 ( .gnd(gnd), .vdd(vdd), .A(_3667__76_), .Y(_1733_) );
OAI21X1 OAI21X1_1070 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1733_), .Y(_1734_) );
AOI22X1 AOI22X1_717 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(b_reg_14_), .C(_1734_), .D(_3433__bF_buf7), .Y(_1735_) );
OAI21X1 OAI21X1_1071 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_3387__bF_buf4), .C(_1735_), .Y(_7__12_) );
INVX1 INVX1_792 ( .gnd(gnd), .vdd(vdd), .A(_3667__77_), .Y(_1736_) );
NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_3432__bF_buf4), .Y(_1737_) );
AOI22X1 AOI22X1_718 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(b_reg_15_), .C(_3433__bF_buf6), .D(_1737_), .Y(_1738_) );
OAI21X1 OAI21X1_1072 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_3387__bF_buf3), .C(_1738_), .Y(_7__13_) );
INVX1 INVX1_793 ( .gnd(gnd), .vdd(vdd), .A(c_reg_14_), .Y(_1739_) );
INVX1 INVX1_794 ( .gnd(gnd), .vdd(vdd), .A(_3667__78_), .Y(_1740_) );
OAI21X1 OAI21X1_1073 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1740_), .Y(_1741_) );
AOI22X1 AOI22X1_719 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(b_reg_16_), .C(_1741_), .D(_3433__bF_buf5), .Y(_1742_) );
OAI21X1 OAI21X1_1074 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_3387__bF_buf2), .C(_1742_), .Y(_7__14_) );
INVX1 INVX1_795 ( .gnd(gnd), .vdd(vdd), .A(_3667__79_), .Y(_1743_) );
OAI21X1 OAI21X1_1075 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1743_), .Y(_1744_) );
AOI22X1 AOI22X1_720 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(b_reg_17_), .C(_1744_), .D(_3433__bF_buf4), .Y(_1745_) );
OAI21X1 OAI21X1_1076 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_3387__bF_buf1), .C(_1745_), .Y(_7__15_) );
INVX1 INVX1_796 ( .gnd(gnd), .vdd(vdd), .A(_3667__80_), .Y(_1746_) );
NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .B(_3432__bF_buf3), .Y(_1747_) );
AOI22X1 AOI22X1_721 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(b_reg_18_), .C(_3433__bF_buf3), .D(_1747_), .Y(_1748_) );
OAI21X1 OAI21X1_1077 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_3387__bF_buf0), .C(_1748_), .Y(_7__16_) );
INVX1 INVX1_797 ( .gnd(gnd), .vdd(vdd), .A(_3667__81_), .Y(_1749_) );
OAI21X1 OAI21X1_1078 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1749_), .Y(_1750_) );
AOI22X1 AOI22X1_722 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(b_reg_19_), .C(_1750_), .D(_3433__bF_buf2), .Y(_1751_) );
OAI21X1 OAI21X1_1079 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_3387__bF_buf10), .C(_1751_), .Y(_7__17_) );
INVX1 INVX1_798 ( .gnd(gnd), .vdd(vdd), .A(_3667__82_), .Y(_1752_) );
NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_3432__bF_buf2), .Y(_1753_) );
AOI22X1 AOI22X1_723 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(b_reg_20_), .C(_3433__bF_buf1), .D(_1753_), .Y(_1754_) );
OAI21X1 OAI21X1_1080 ( .gnd(gnd), .vdd(vdd), .A(_908_), .B(_3387__bF_buf9), .C(_1754_), .Y(_7__18_) );
INVX1 INVX1_799 ( .gnd(gnd), .vdd(vdd), .A(_3667__83_), .Y(_1755_) );
OAI21X1 OAI21X1_1081 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1755_), .Y(_1756_) );
AOI22X1 AOI22X1_724 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(b_reg_21_), .C(_1756_), .D(_3433__bF_buf0), .Y(_1757_) );
OAI21X1 OAI21X1_1082 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_3387__bF_buf8), .C(_1757_), .Y(_7__19_) );
INVX1 INVX1_800 ( .gnd(gnd), .vdd(vdd), .A(_3667__84_), .Y(_1758_) );
OAI21X1 OAI21X1_1083 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1758_), .Y(_1759_) );
AOI22X1 AOI22X1_725 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(b_reg_22_), .C(_1759_), .D(_3433__bF_buf11), .Y(_1760_) );
OAI21X1 OAI21X1_1084 ( .gnd(gnd), .vdd(vdd), .A(_1022_), .B(_3387__bF_buf7), .C(_1760_), .Y(_7__20_) );
INVX1 INVX1_801 ( .gnd(gnd), .vdd(vdd), .A(_3667__85_), .Y(_1761_) );
OAI21X1 OAI21X1_1085 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1761_), .Y(_1762_) );
AOI22X1 AOI22X1_726 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(b_reg_23_), .C(_1762_), .D(_3433__bF_buf10), .Y(_1763_) );
OAI21X1 OAI21X1_1086 ( .gnd(gnd), .vdd(vdd), .A(_1082_), .B(_3387__bF_buf6), .C(_1763_), .Y(_7__21_) );
INVX1 INVX1_802 ( .gnd(gnd), .vdd(vdd), .A(_3667__86_), .Y(_1764_) );
NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(_1764_), .B(_3432__bF_buf1), .Y(_1765_) );
AOI22X1 AOI22X1_727 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(b_reg_24_), .C(_3433__bF_buf9), .D(_1765_), .Y(_1766_) );
OAI21X1 OAI21X1_1087 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_3387__bF_buf5), .C(_1766_), .Y(_7__22_) );
INVX1 INVX1_803 ( .gnd(gnd), .vdd(vdd), .A(_3667__87_), .Y(_1767_) );
OAI21X1 OAI21X1_1088 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1767_), .Y(_1769_) );
AOI22X1 AOI22X1_728 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(b_reg_25_), .C(_1769_), .D(_3433__bF_buf8), .Y(_1770_) );
OAI21X1 OAI21X1_1089 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_3387__bF_buf4), .C(_1770_), .Y(_7__23_) );
INVX1 INVX1_804 ( .gnd(gnd), .vdd(vdd), .A(_3667__88_), .Y(_1771_) );
NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .B(_3432__bF_buf0), .Y(_1772_) );
AOI22X1 AOI22X1_729 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(b_reg_26_), .C(_3433__bF_buf7), .D(_1772_), .Y(_1773_) );
OAI21X1 OAI21X1_1090 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_3387__bF_buf3), .C(_1773_), .Y(_7__24_) );
INVX1 INVX1_805 ( .gnd(gnd), .vdd(vdd), .A(_3667__89_), .Y(_1774_) );
NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_3432__bF_buf11), .Y(_1775_) );
AOI22X1 AOI22X1_730 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(b_reg_27_), .C(_3433__bF_buf6), .D(_1775_), .Y(_1776_) );
OAI21X1 OAI21X1_1091 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_3387__bF_buf2), .C(_1776_), .Y(_7__25_) );
INVX2 INVX2_72 ( .gnd(gnd), .vdd(vdd), .A(_3667__90_), .Y(_1777_) );
NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_3432__bF_buf10), .Y(_1778_) );
AOI22X1 AOI22X1_731 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(b_reg_28_), .C(_3433__bF_buf5), .D(_1778_), .Y(_1779_) );
OAI21X1 OAI21X1_1092 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_3387__bF_buf1), .C(_1779_), .Y(_7__26_) );
INVX1 INVX1_806 ( .gnd(gnd), .vdd(vdd), .A(_3667__91_), .Y(_1780_) );
OAI21X1 OAI21X1_1093 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1780_), .Y(_1781_) );
AOI22X1 AOI22X1_732 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(b_reg_29_), .C(_1781_), .D(_3433__bF_buf4), .Y(_1782_) );
OAI21X1 OAI21X1_1094 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_3387__bF_buf0), .C(_1782_), .Y(_7__27_) );
INVX1 INVX1_807 ( .gnd(gnd), .vdd(vdd), .A(_3667__92_), .Y(_1783_) );
OAI21X1 OAI21X1_1095 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1783_), .Y(_1784_) );
AOI22X1 AOI22X1_733 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(b_reg_30_), .C(_1784_), .D(_3433__bF_buf3), .Y(_1785_) );
OAI21X1 OAI21X1_1096 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_3387__bF_buf10), .C(_1785_), .Y(_7__28_) );
INVX1 INVX1_808 ( .gnd(gnd), .vdd(vdd), .A(_3667__93_), .Y(_1786_) );
NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(_1786_), .B(_3432__bF_buf9), .Y(_1787_) );
AOI22X1 AOI22X1_734 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(b_reg_31_), .C(_3433__bF_buf2), .D(_1787_), .Y(_1788_) );
OAI21X1 OAI21X1_1097 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(_3387__bF_buf9), .C(_1788_), .Y(_7__29_) );
INVX2 INVX2_73 ( .gnd(gnd), .vdd(vdd), .A(_3667__94_), .Y(_1789_) );
NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_3432__bF_buf8), .Y(_1790_) );
AOI22X1 AOI22X1_735 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(b_reg_0_), .C(_3433__bF_buf1), .D(_1790_), .Y(_1791_) );
OAI21X1 OAI21X1_1098 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_3387__bF_buf8), .C(_1791_), .Y(_7__30_) );
OAI21X1 OAI21X1_1099 ( .gnd(gnd), .vdd(vdd), .A(_3667__95_), .B(_3432__bF_buf7), .C(_3433__bF_buf0), .Y(_1792_) );
AOI22X1 AOI22X1_736 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(b_reg_1_), .C(c_reg_31_), .D(_113__bF_buf2), .Y(_1793_) );
NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_1792_), .B(_1793_), .Y(_7__31_) );
INVX1 INVX1_809 ( .gnd(gnd), .vdd(vdd), .A(_3667__32_), .Y(_1794_) );
NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(_3432__bF_buf6), .Y(_1795_) );
AOI22X1 AOI22X1_737 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(c_reg_0_), .C(_3433__bF_buf11), .D(_1795_), .Y(_1796_) );
OAI21X1 OAI21X1_1100 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_3387__bF_buf7), .C(_1796_), .Y(_8__0_) );
INVX1 INVX1_810 ( .gnd(gnd), .vdd(vdd), .A(_3667__33_), .Y(_1797_) );
OAI21X1 OAI21X1_1101 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1797_), .Y(_1798_) );
AOI22X1 AOI22X1_738 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(c_reg_1_), .C(_1798_), .D(_3433__bF_buf10), .Y(_1799_) );
OAI21X1 OAI21X1_1102 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_3387__bF_buf6), .C(_1799_), .Y(_8__1_) );
INVX1 INVX1_811 ( .gnd(gnd), .vdd(vdd), .A(_3667__34_), .Y(_1800_) );
OAI21X1 OAI21X1_1103 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1800_), .Y(_1801_) );
AOI22X1 AOI22X1_739 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(c_reg_2_), .C(_1801_), .D(_3433__bF_buf9), .Y(_1802_) );
OAI21X1 OAI21X1_1104 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_3387__bF_buf5), .C(_1802_), .Y(_8__2_) );
INVX1 INVX1_812 ( .gnd(gnd), .vdd(vdd), .A(_3667__35_), .Y(_1803_) );
NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_3432__bF_buf5), .Y(_1804_) );
AOI22X1 AOI22X1_740 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(c_reg_3_), .C(_3433__bF_buf8), .D(_1804_), .Y(_1805_) );
OAI21X1 OAI21X1_1105 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_3387__bF_buf4), .C(_1805_), .Y(_8__3_) );
INVX1 INVX1_813 ( .gnd(gnd), .vdd(vdd), .A(_3667__36_), .Y(_1806_) );
OAI21X1 OAI21X1_1106 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1806_), .Y(_1807_) );
AOI22X1 AOI22X1_741 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(c_reg_4_), .C(_1807_), .D(_3433__bF_buf7), .Y(_1808_) );
OAI21X1 OAI21X1_1107 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(_3387__bF_buf3), .C(_1808_), .Y(_8__4_) );
INVX1 INVX1_814 ( .gnd(gnd), .vdd(vdd), .A(_3667__37_), .Y(_1809_) );
OAI21X1 OAI21X1_1108 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1809_), .Y(_1810_) );
AOI22X1 AOI22X1_742 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(c_reg_5_), .C(_1810_), .D(_3433__bF_buf6), .Y(_1811_) );
OAI21X1 OAI21X1_1109 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_3387__bF_buf2), .C(_1811_), .Y(_8__5_) );
INVX1 INVX1_815 ( .gnd(gnd), .vdd(vdd), .A(_3667__38_), .Y(_1812_) );
OAI21X1 OAI21X1_1110 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1812_), .Y(_1813_) );
AOI22X1 AOI22X1_743 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(c_reg_6_), .C(_1813_), .D(_3433__bF_buf5), .Y(_1814_) );
OAI21X1 OAI21X1_1111 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_3387__bF_buf1), .C(_1814_), .Y(_8__6_) );
INVX1 INVX1_816 ( .gnd(gnd), .vdd(vdd), .A(_3667__39_), .Y(_1815_) );
NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(_3432__bF_buf4), .Y(_1816_) );
AOI22X1 AOI22X1_744 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(c_reg_7_), .C(_3433__bF_buf4), .D(_1816_), .Y(_1817_) );
OAI21X1 OAI21X1_1112 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_3387__bF_buf0), .C(_1817_), .Y(_8__7_) );
INVX1 INVX1_817 ( .gnd(gnd), .vdd(vdd), .A(_3667__40_), .Y(_1818_) );
NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_3432__bF_buf3), .Y(_1819_) );
AOI22X1 AOI22X1_745 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(c_reg_8_), .C(_3433__bF_buf3), .D(_1819_), .Y(_1820_) );
OAI21X1 OAI21X1_1113 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_3387__bF_buf10), .C(_1820_), .Y(_8__8_) );
INVX1 INVX1_818 ( .gnd(gnd), .vdd(vdd), .A(_3667__41_), .Y(_1821_) );
NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_3432__bF_buf2), .Y(_1822_) );
AOI22X1 AOI22X1_746 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(c_reg_9_), .C(_3433__bF_buf2), .D(_1822_), .Y(_1823_) );
OAI21X1 OAI21X1_1114 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_3387__bF_buf9), .C(_1823_), .Y(_8__9_) );
INVX1 INVX1_819 ( .gnd(gnd), .vdd(vdd), .A(_3667__42_), .Y(_1824_) );
OAI21X1 OAI21X1_1115 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1824_), .Y(_1825_) );
AOI22X1 AOI22X1_747 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(c_reg_10_), .C(_1825_), .D(_3433__bF_buf1), .Y(_1826_) );
OAI21X1 OAI21X1_1116 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_3387__bF_buf8), .C(_1826_), .Y(_8__10_) );
INVX1 INVX1_820 ( .gnd(gnd), .vdd(vdd), .A(_3667__43_), .Y(_1827_) );
NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_3432__bF_buf1), .Y(_1828_) );
AOI22X1 AOI22X1_748 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(c_reg_11_), .C(_3433__bF_buf0), .D(_1828_), .Y(_1829_) );
OAI21X1 OAI21X1_1117 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_3387__bF_buf7), .C(_1829_), .Y(_8__11_) );
INVX1 INVX1_821 ( .gnd(gnd), .vdd(vdd), .A(_3667__44_), .Y(_1830_) );
OAI21X1 OAI21X1_1118 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1830_), .Y(_1831_) );
AOI22X1 AOI22X1_749 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(c_reg_12_), .C(_1831_), .D(_3433__bF_buf11), .Y(_1832_) );
OAI21X1 OAI21X1_1119 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_3387__bF_buf6), .C(_1832_), .Y(_8__12_) );
INVX2 INVX2_74 ( .gnd(gnd), .vdd(vdd), .A(_3667__45_), .Y(_1833_) );
NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_3432__bF_buf0), .Y(_1834_) );
AOI22X1 AOI22X1_750 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(c_reg_13_), .C(_3433__bF_buf10), .D(_1834_), .Y(_1835_) );
OAI21X1 OAI21X1_1120 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_3387__bF_buf5), .C(_1835_), .Y(_8__13_) );
INVX1 INVX1_822 ( .gnd(gnd), .vdd(vdd), .A(_3667__46_), .Y(_1836_) );
OAI21X1 OAI21X1_1121 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1836_), .Y(_1837_) );
AOI22X1 AOI22X1_751 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(c_reg_14_), .C(_1837_), .D(_3433__bF_buf9), .Y(_1838_) );
OAI21X1 OAI21X1_1122 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_3387__bF_buf4), .C(_1838_), .Y(_8__14_) );
INVX1 INVX1_823 ( .gnd(gnd), .vdd(vdd), .A(_3667__47_), .Y(_1839_) );
NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_3432__bF_buf11), .Y(_1840_) );
AOI22X1 AOI22X1_752 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(c_reg_15_), .C(_3433__bF_buf8), .D(_1840_), .Y(_1841_) );
OAI21X1 OAI21X1_1123 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_3387__bF_buf3), .C(_1841_), .Y(_8__15_) );
INVX1 INVX1_824 ( .gnd(gnd), .vdd(vdd), .A(_3667__48_), .Y(_1842_) );
NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_3432__bF_buf10), .Y(_1843_) );
AOI22X1 AOI22X1_753 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(c_reg_16_), .C(_3433__bF_buf7), .D(_1843_), .Y(_1844_) );
OAI21X1 OAI21X1_1124 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_3387__bF_buf2), .C(_1844_), .Y(_8__16_) );
INVX1 INVX1_825 ( .gnd(gnd), .vdd(vdd), .A(_3667__49_), .Y(_1845_) );
OAI21X1 OAI21X1_1125 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1845_), .Y(_1846_) );
AOI22X1 AOI22X1_754 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(c_reg_17_), .C(_1846_), .D(_3433__bF_buf6), .Y(_1847_) );
OAI21X1 OAI21X1_1126 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_3387__bF_buf1), .C(_1847_), .Y(_8__17_) );
INVX1 INVX1_826 ( .gnd(gnd), .vdd(vdd), .A(_3667__50_), .Y(_1848_) );
NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_3432__bF_buf9), .Y(_1849_) );
AOI22X1 AOI22X1_755 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(c_reg_18_), .C(_3433__bF_buf5), .D(_1849_), .Y(_1850_) );
OAI21X1 OAI21X1_1127 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_3387__bF_buf0), .C(_1850_), .Y(_8__18_) );
INVX1 INVX1_827 ( .gnd(gnd), .vdd(vdd), .A(_3667__51_), .Y(_1851_) );
NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(_3432__bF_buf8), .Y(_1852_) );
AOI22X1 AOI22X1_756 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(c_reg_19_), .C(_3433__bF_buf4), .D(_1852_), .Y(_1853_) );
OAI21X1 OAI21X1_1128 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_3387__bF_buf10), .C(_1853_), .Y(_8__19_) );
INVX1 INVX1_828 ( .gnd(gnd), .vdd(vdd), .A(_3667__52_), .Y(_1854_) );
OAI21X1 OAI21X1_1129 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1854_), .Y(_1855_) );
AOI22X1 AOI22X1_757 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(c_reg_20_), .C(_1855_), .D(_3433__bF_buf3), .Y(_1856_) );
OAI21X1 OAI21X1_1130 ( .gnd(gnd), .vdd(vdd), .A(_1024_), .B(_3387__bF_buf9), .C(_1856_), .Y(_8__20_) );
INVX1 INVX1_829 ( .gnd(gnd), .vdd(vdd), .A(_3667__53_), .Y(_1857_) );
OAI21X1 OAI21X1_1131 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1857_), .Y(_1858_) );
AOI22X1 AOI22X1_758 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(c_reg_21_), .C(_1858_), .D(_3433__bF_buf2), .Y(_1859_) );
OAI21X1 OAI21X1_1132 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_3387__bF_buf8), .C(_1859_), .Y(_8__21_) );
INVX1 INVX1_830 ( .gnd(gnd), .vdd(vdd), .A(_3667__54_), .Y(_1860_) );
NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_3432__bF_buf7), .Y(_1861_) );
AOI22X1 AOI22X1_759 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(c_reg_22_), .C(_3433__bF_buf1), .D(_1861_), .Y(_1862_) );
OAI21X1 OAI21X1_1133 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(_3387__bF_buf7), .C(_1862_), .Y(_8__22_) );
INVX1 INVX1_831 ( .gnd(gnd), .vdd(vdd), .A(_3667__55_), .Y(_1863_) );
NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_3432__bF_buf6), .Y(_1864_) );
AOI22X1 AOI22X1_760 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(c_reg_23_), .C(_3433__bF_buf0), .D(_1864_), .Y(_1865_) );
OAI21X1 OAI21X1_1134 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_3387__bF_buf6), .C(_1865_), .Y(_8__23_) );
INVX1 INVX1_832 ( .gnd(gnd), .vdd(vdd), .A(_3667__56_), .Y(_1866_) );
NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(_3432__bF_buf5), .Y(_1867_) );
AOI22X1 AOI22X1_761 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(c_reg_24_), .C(_3433__bF_buf11), .D(_1867_), .Y(_1868_) );
OAI21X1 OAI21X1_1135 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_3387__bF_buf5), .C(_1868_), .Y(_8__24_) );
INVX2 INVX2_75 ( .gnd(gnd), .vdd(vdd), .A(_3667__57_), .Y(_1869_) );
NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(_1869_), .B(_3432__bF_buf4), .Y(_1870_) );
AOI22X1 AOI22X1_762 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(c_reg_25_), .C(_3433__bF_buf10), .D(_1870_), .Y(_1871_) );
OAI21X1 OAI21X1_1136 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_3387__bF_buf4), .C(_1871_), .Y(_8__25_) );
INVX1 INVX1_833 ( .gnd(gnd), .vdd(vdd), .A(_3667__58_), .Y(_1872_) );
NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(_1872_), .B(_3432__bF_buf3), .Y(_1873_) );
AOI22X1 AOI22X1_763 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(c_reg_26_), .C(_3433__bF_buf9), .D(_1873_), .Y(_1874_) );
OAI21X1 OAI21X1_1137 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_3387__bF_buf3), .C(_1874_), .Y(_8__26_) );
INVX1 INVX1_834 ( .gnd(gnd), .vdd(vdd), .A(d_reg_27_), .Y(_1875_) );
INVX2 INVX2_76 ( .gnd(gnd), .vdd(vdd), .A(_3667__59_), .Y(_1876_) );
NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(_1876_), .B(_3432__bF_buf2), .Y(_1877_) );
AOI22X1 AOI22X1_764 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(c_reg_27_), .C(_3433__bF_buf8), .D(_1877_), .Y(_1878_) );
OAI21X1 OAI21X1_1138 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(_3387__bF_buf2), .C(_1878_), .Y(_8__27_) );
INVX1 INVX1_835 ( .gnd(gnd), .vdd(vdd), .A(_3667__60_), .Y(_1879_) );
OAI21X1 OAI21X1_1139 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1879_), .Y(_1880_) );
AOI22X1 AOI22X1_765 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(c_reg_28_), .C(_1880_), .D(_3433__bF_buf7), .Y(_1881_) );
OAI21X1 OAI21X1_1140 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_3387__bF_buf1), .C(_1881_), .Y(_8__28_) );
INVX1 INVX1_836 ( .gnd(gnd), .vdd(vdd), .A(_3667__61_), .Y(_1882_) );
NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(_1882_), .B(_3432__bF_buf1), .Y(_1883_) );
AOI22X1 AOI22X1_766 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(c_reg_29_), .C(_3433__bF_buf6), .D(_1883_), .Y(_1884_) );
OAI21X1 OAI21X1_1141 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_3387__bF_buf0), .C(_1884_), .Y(_8__29_) );
INVX2 INVX2_77 ( .gnd(gnd), .vdd(vdd), .A(_3667__62_), .Y(_1885_) );
NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(_1885_), .B(_3432__bF_buf0), .Y(_1886_) );
AOI22X1 AOI22X1_767 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(c_reg_30_), .C(_3433__bF_buf5), .D(_1886_), .Y(_1887_) );
OAI21X1 OAI21X1_1142 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_3387__bF_buf10), .C(_1887_), .Y(_8__30_) );
INVX1 INVX1_837 ( .gnd(gnd), .vdd(vdd), .A(_3432__bF_buf11), .Y(_1888_) );
NAND3X1 NAND3X1_291 ( .gnd(gnd), .vdd(vdd), .A(_3667__63_), .B(_3433__bF_buf4), .C(_1888_), .Y(_1889_) );
NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(d_reg_31_), .B(_113__bF_buf1), .Y(_1890_) );
NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(c_reg_31_), .Y(_1891_) );
NAND3X1 NAND3X1_292 ( .gnd(gnd), .vdd(vdd), .A(_1891_), .B(_1889_), .C(_1890_), .Y(_8__31_) );
INVX1 INVX1_838 ( .gnd(gnd), .vdd(vdd), .A(e_reg_0_), .Y(_1892_) );
INVX1 INVX1_839 ( .gnd(gnd), .vdd(vdd), .A(_3667__0_), .Y(_1893_) );
NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(_1893_), .B(_3432__bF_buf10), .Y(_1894_) );
AOI22X1 AOI22X1_768 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(d_reg_0_), .C(_3433__bF_buf3), .D(_1894_), .Y(_1895_) );
OAI21X1 OAI21X1_1143 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_3387__bF_buf9), .C(_1895_), .Y(_10__0_) );
INVX1 INVX1_840 ( .gnd(gnd), .vdd(vdd), .A(e_reg_1_), .Y(_1896_) );
INVX1 INVX1_841 ( .gnd(gnd), .vdd(vdd), .A(_3667__1_), .Y(_1897_) );
NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(_3432__bF_buf9), .Y(_1898_) );
AOI22X1 AOI22X1_769 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(d_reg_1_), .C(_3433__bF_buf2), .D(_1898_), .Y(_1899_) );
OAI21X1 OAI21X1_1144 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(_3387__bF_buf8), .C(_1899_), .Y(_10__1_) );
INVX1 INVX1_842 ( .gnd(gnd), .vdd(vdd), .A(e_reg_2_), .Y(_1900_) );
INVX1 INVX1_843 ( .gnd(gnd), .vdd(vdd), .A(_3667__2_), .Y(_1901_) );
NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .B(_3432__bF_buf8), .Y(_1902_) );
AOI22X1 AOI22X1_770 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(d_reg_2_), .C(_3433__bF_buf1), .D(_1902_), .Y(_1903_) );
OAI21X1 OAI21X1_1145 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(_3387__bF_buf7), .C(_1903_), .Y(_10__2_) );
INVX1 INVX1_844 ( .gnd(gnd), .vdd(vdd), .A(e_reg_3_), .Y(_1904_) );
INVX1 INVX1_845 ( .gnd(gnd), .vdd(vdd), .A(_3667__3_), .Y(_1905_) );
NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(_3432__bF_buf7), .Y(_1906_) );
AOI22X1 AOI22X1_771 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(d_reg_3_), .C(_3433__bF_buf0), .D(_1906_), .Y(_1907_) );
OAI21X1 OAI21X1_1146 ( .gnd(gnd), .vdd(vdd), .A(_1904_), .B(_3387__bF_buf6), .C(_1907_), .Y(_10__3_) );
INVX1 INVX1_846 ( .gnd(gnd), .vdd(vdd), .A(e_reg_4_), .Y(_1908_) );
INVX1 INVX1_847 ( .gnd(gnd), .vdd(vdd), .A(_3667__4_), .Y(_1909_) );
OAI21X1 OAI21X1_1147 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1909_), .Y(_1910_) );
AOI22X1 AOI22X1_772 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(d_reg_4_), .C(_1910_), .D(_3433__bF_buf11), .Y(_1911_) );
OAI21X1 OAI21X1_1148 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(_3387__bF_buf5), .C(_1911_), .Y(_10__4_) );
INVX1 INVX1_848 ( .gnd(gnd), .vdd(vdd), .A(_3667__5_), .Y(_1912_) );
OAI21X1 OAI21X1_1149 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1912_), .Y(_1913_) );
AOI22X1 AOI22X1_773 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(d_reg_5_), .C(_1913_), .D(_3433__bF_buf10), .Y(_1914_) );
OAI21X1 OAI21X1_1150 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_3387__bF_buf4), .C(_1914_), .Y(_10__5_) );
INVX1 INVX1_849 ( .gnd(gnd), .vdd(vdd), .A(e_reg_6_), .Y(_1915_) );
INVX1 INVX1_850 ( .gnd(gnd), .vdd(vdd), .A(_3667__6_), .Y(_1916_) );
OAI21X1 OAI21X1_1151 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1916_), .Y(_1917_) );
AOI22X1 AOI22X1_774 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(d_reg_6_), .C(_1917_), .D(_3433__bF_buf9), .Y(_1918_) );
OAI21X1 OAI21X1_1152 ( .gnd(gnd), .vdd(vdd), .A(_1915_), .B(_3387__bF_buf3), .C(_1918_), .Y(_10__6_) );
OAI21X1 OAI21X1_1153 ( .gnd(gnd), .vdd(vdd), .A(_3667__7_), .B(_3432__bF_buf6), .C(_3433__bF_buf8), .Y(_1919_) );
AOI22X1 AOI22X1_775 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(d_reg_7_), .C(e_reg_7_), .D(_113__bF_buf0), .Y(_1920_) );
NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(_1919_), .B(_1920_), .Y(_10__7_) );
INVX1 INVX1_851 ( .gnd(gnd), .vdd(vdd), .A(e_reg_8_), .Y(_1921_) );
INVX1 INVX1_852 ( .gnd(gnd), .vdd(vdd), .A(_3667__8_), .Y(_1922_) );
OAI21X1 OAI21X1_1154 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1922_), .Y(_1923_) );
AOI22X1 AOI22X1_776 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(d_reg_8_), .C(_1923_), .D(_3433__bF_buf7), .Y(_1924_) );
OAI21X1 OAI21X1_1155 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_3387__bF_buf2), .C(_1924_), .Y(_10__8_) );
INVX1 INVX1_853 ( .gnd(gnd), .vdd(vdd), .A(e_reg_9_), .Y(_1925_) );
INVX2 INVX2_78 ( .gnd(gnd), .vdd(vdd), .A(_3667__9_), .Y(_1926_) );
NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_3432__bF_buf5), .Y(_1927_) );
AOI22X1 AOI22X1_777 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(d_reg_9_), .C(_3433__bF_buf6), .D(_1927_), .Y(_1928_) );
OAI21X1 OAI21X1_1156 ( .gnd(gnd), .vdd(vdd), .A(_1925_), .B(_3387__bF_buf1), .C(_1928_), .Y(_10__9_) );
INVX1 INVX1_854 ( .gnd(gnd), .vdd(vdd), .A(e_reg_10_), .Y(_1929_) );
INVX1 INVX1_855 ( .gnd(gnd), .vdd(vdd), .A(_3667__10_), .Y(_1930_) );
NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_3432__bF_buf4), .Y(_1931_) );
AOI22X1 AOI22X1_778 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(d_reg_10_), .C(_3433__bF_buf5), .D(_1931_), .Y(_1932_) );
OAI21X1 OAI21X1_1157 ( .gnd(gnd), .vdd(vdd), .A(_1929_), .B(_3387__bF_buf0), .C(_1932_), .Y(_10__10_) );
INVX1 INVX1_856 ( .gnd(gnd), .vdd(vdd), .A(e_reg_11_), .Y(_1933_) );
INVX1 INVX1_857 ( .gnd(gnd), .vdd(vdd), .A(_3667__11_), .Y(_1934_) );
NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .B(_3432__bF_buf3), .Y(_1935_) );
AOI22X1 AOI22X1_779 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(d_reg_11_), .C(_3433__bF_buf4), .D(_1935_), .Y(_1936_) );
OAI21X1 OAI21X1_1158 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .B(_3387__bF_buf10), .C(_1936_), .Y(_10__11_) );
INVX1 INVX1_858 ( .gnd(gnd), .vdd(vdd), .A(e_reg_12_), .Y(_1937_) );
INVX2 INVX2_79 ( .gnd(gnd), .vdd(vdd), .A(_3667__12_), .Y(_1938_) );
NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_3432__bF_buf2), .Y(_1939_) );
AOI22X1 AOI22X1_780 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(d_reg_12_), .C(_3433__bF_buf3), .D(_1939_), .Y(_1940_) );
OAI21X1 OAI21X1_1159 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .B(_3387__bF_buf9), .C(_1940_), .Y(_10__12_) );
INVX1 INVX1_859 ( .gnd(gnd), .vdd(vdd), .A(e_reg_13_), .Y(_1941_) );
INVX1 INVX1_860 ( .gnd(gnd), .vdd(vdd), .A(_3667__13_), .Y(_1942_) );
OAI21X1 OAI21X1_1160 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1942_), .Y(_1943_) );
AOI22X1 AOI22X1_781 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(d_reg_13_), .C(_1943_), .D(_3433__bF_buf2), .Y(_1944_) );
OAI21X1 OAI21X1_1161 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(_3387__bF_buf8), .C(_1944_), .Y(_10__13_) );
INVX1 INVX1_861 ( .gnd(gnd), .vdd(vdd), .A(e_reg_14_), .Y(_1945_) );
INVX1 INVX1_862 ( .gnd(gnd), .vdd(vdd), .A(_3667__14_), .Y(_1946_) );
OAI21X1 OAI21X1_1162 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_1946_), .Y(_1947_) );
AOI22X1 AOI22X1_782 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(d_reg_14_), .C(_1947_), .D(_3433__bF_buf1), .Y(_1948_) );
OAI21X1 OAI21X1_1163 ( .gnd(gnd), .vdd(vdd), .A(_1945_), .B(_3387__bF_buf7), .C(_1948_), .Y(_10__14_) );
INVX1 INVX1_863 ( .gnd(gnd), .vdd(vdd), .A(e_reg_15_), .Y(_1949_) );
INVX1 INVX1_864 ( .gnd(gnd), .vdd(vdd), .A(_3667__15_), .Y(_1950_) );
OAI21X1 OAI21X1_1164 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf1), .B(_3386__bF_buf0), .C(_1950_), .Y(_1951_) );
AOI22X1 AOI22X1_783 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(d_reg_15_), .C(_1951_), .D(_3433__bF_buf0), .Y(_1952_) );
OAI21X1 OAI21X1_1165 ( .gnd(gnd), .vdd(vdd), .A(_1949_), .B(_3387__bF_buf6), .C(_1952_), .Y(_10__15_) );
INVX1 INVX1_865 ( .gnd(gnd), .vdd(vdd), .A(_3667__16_), .Y(_1953_) );
NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(_1953_), .B(_3432__bF_buf1), .Y(_1954_) );
AOI22X1 AOI22X1_784 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(d_reg_16_), .C(_3433__bF_buf11), .D(_1954_), .Y(_1955_) );
OAI21X1 OAI21X1_1166 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_3387__bF_buf5), .C(_1955_), .Y(_10__16_) );
INVX1 INVX1_866 ( .gnd(gnd), .vdd(vdd), .A(e_reg_17_), .Y(_1956_) );
INVX1 INVX1_867 ( .gnd(gnd), .vdd(vdd), .A(_3667__17_), .Y(_1957_) );
OAI21X1 OAI21X1_1167 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf0), .B(_3386__bF_buf7), .C(_1957_), .Y(_1958_) );
AOI22X1 AOI22X1_785 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(d_reg_17_), .C(_1958_), .D(_3433__bF_buf10), .Y(_1959_) );
OAI21X1 OAI21X1_1168 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_3387__bF_buf4), .C(_1959_), .Y(_10__17_) );
INVX1 INVX1_868 ( .gnd(gnd), .vdd(vdd), .A(_3667__18_), .Y(_1960_) );
NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .B(_3432__bF_buf0), .Y(_1961_) );
AOI22X1 AOI22X1_786 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(d_reg_18_), .C(_3433__bF_buf9), .D(_1961_), .Y(_1962_) );
OAI21X1 OAI21X1_1169 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_3387__bF_buf3), .C(_1962_), .Y(_10__18_) );
INVX1 INVX1_869 ( .gnd(gnd), .vdd(vdd), .A(e_reg_19_), .Y(_1963_) );
INVX1 INVX1_870 ( .gnd(gnd), .vdd(vdd), .A(_3667__19_), .Y(_1964_) );
NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(_3432__bF_buf11), .Y(_1965_) );
AOI22X1 AOI22X1_787 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(d_reg_19_), .C(_3433__bF_buf8), .D(_1965_), .Y(_1966_) );
OAI21X1 OAI21X1_1170 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_3387__bF_buf2), .C(_1966_), .Y(_10__19_) );
INVX1 INVX1_871 ( .gnd(gnd), .vdd(vdd), .A(e_reg_20_), .Y(_1967_) );
INVX1 INVX1_872 ( .gnd(gnd), .vdd(vdd), .A(_3667__20_), .Y(_1968_) );
OAI21X1 OAI21X1_1171 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf7), .B(_3386__bF_buf6), .C(_1968_), .Y(_1969_) );
AOI22X1 AOI22X1_788 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(d_reg_20_), .C(_1969_), .D(_3433__bF_buf7), .Y(_1970_) );
OAI21X1 OAI21X1_1172 ( .gnd(gnd), .vdd(vdd), .A(_1967_), .B(_3387__bF_buf1), .C(_1970_), .Y(_10__20_) );
INVX1 INVX1_873 ( .gnd(gnd), .vdd(vdd), .A(e_reg_21_), .Y(_1971_) );
INVX2 INVX2_80 ( .gnd(gnd), .vdd(vdd), .A(_3667__21_), .Y(_1972_) );
NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(_1972_), .B(_3432__bF_buf10), .Y(_1973_) );
AOI22X1 AOI22X1_789 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(d_reg_21_), .C(_3433__bF_buf6), .D(_1973_), .Y(_1974_) );
OAI21X1 OAI21X1_1173 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_3387__bF_buf0), .C(_1974_), .Y(_10__21_) );
INVX1 INVX1_874 ( .gnd(gnd), .vdd(vdd), .A(_3667__22_), .Y(_1975_) );
OAI21X1 OAI21X1_1174 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf6), .B(_3386__bF_buf5), .C(_1975_), .Y(_1976_) );
AOI22X1 AOI22X1_790 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(d_reg_22_), .C(_1976_), .D(_3433__bF_buf5), .Y(_1977_) );
OAI21X1 OAI21X1_1175 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_3387__bF_buf10), .C(_1977_), .Y(_10__22_) );
INVX1 INVX1_875 ( .gnd(gnd), .vdd(vdd), .A(_3667__23_), .Y(_1978_) );
OAI21X1 OAI21X1_1176 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf5), .B(_3386__bF_buf4), .C(_1978_), .Y(_1979_) );
AOI22X1 AOI22X1_791 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(d_reg_23_), .C(_1979_), .D(_3433__bF_buf4), .Y(_1980_) );
OAI21X1 OAI21X1_1177 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_3387__bF_buf9), .C(_1980_), .Y(_10__23_) );
INVX1 INVX1_876 ( .gnd(gnd), .vdd(vdd), .A(_3667__24_), .Y(_1981_) );
OAI21X1 OAI21X1_1178 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf4), .B(_3386__bF_buf3), .C(_1981_), .Y(_1982_) );
AOI22X1 AOI22X1_792 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(d_reg_24_), .C(_1982_), .D(_3433__bF_buf3), .Y(_1983_) );
OAI21X1 OAI21X1_1179 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_3387__bF_buf8), .C(_1983_), .Y(_10__24_) );
INVX1 INVX1_877 ( .gnd(gnd), .vdd(vdd), .A(_3667__25_), .Y(_1984_) );
OAI21X1 OAI21X1_1180 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf3), .B(_3386__bF_buf2), .C(_1984_), .Y(_1985_) );
AOI22X1 AOI22X1_793 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(d_reg_25_), .C(_1985_), .D(_3433__bF_buf2), .Y(_1986_) );
OAI21X1 OAI21X1_1181 ( .gnd(gnd), .vdd(vdd), .A(_1359_), .B(_3387__bF_buf7), .C(_1986_), .Y(_10__25_) );
INVX1 INVX1_878 ( .gnd(gnd), .vdd(vdd), .A(_3667__26_), .Y(_1987_) );
NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(_1987_), .B(_3432__bF_buf9), .Y(_1988_) );
AOI22X1 AOI22X1_794 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf8), .B(d_reg_26_), .C(_3433__bF_buf1), .D(_1988_), .Y(_1989_) );
OAI21X1 OAI21X1_1182 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_3387__bF_buf6), .C(_1989_), .Y(_10__26_) );
INVX1 INVX1_879 ( .gnd(gnd), .vdd(vdd), .A(_3667__27_), .Y(_1990_) );
NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_3432__bF_buf8), .Y(_1991_) );
AOI22X1 AOI22X1_795 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf7), .B(d_reg_27_), .C(_3433__bF_buf0), .D(_1991_), .Y(_1992_) );
OAI21X1 OAI21X1_1183 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_3387__bF_buf5), .C(_1992_), .Y(_10__27_) );
INVX2 INVX2_81 ( .gnd(gnd), .vdd(vdd), .A(_3667__28_), .Y(_1993_) );
NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(_1993_), .B(_3432__bF_buf7), .Y(_1994_) );
AOI22X1 AOI22X1_796 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf6), .B(d_reg_28_), .C(_3433__bF_buf11), .D(_1994_), .Y(_1995_) );
OAI21X1 OAI21X1_1184 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .B(_3387__bF_buf4), .C(_1995_), .Y(_10__28_) );
INVX2 INVX2_82 ( .gnd(gnd), .vdd(vdd), .A(_3667__29_), .Y(_1996_) );
NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_3432__bF_buf6), .Y(_1997_) );
AOI22X1 AOI22X1_797 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf5), .B(d_reg_29_), .C(_3433__bF_buf10), .D(_1997_), .Y(_1998_) );
OAI21X1 OAI21X1_1185 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_3387__bF_buf3), .C(_1998_), .Y(_10__29_) );
OAI21X1 OAI21X1_1186 ( .gnd(gnd), .vdd(vdd), .A(_3667__30_), .B(_3432__bF_buf5), .C(_3433__bF_buf9), .Y(_1999_) );
AOI22X1 AOI22X1_798 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf4), .B(d_reg_30_), .C(e_reg_30_), .D(_113__bF_buf4), .Y(_2000_) );
NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_1999_), .B(_2000_), .Y(_10__30_) );
OAI21X1 OAI21X1_1187 ( .gnd(gnd), .vdd(vdd), .A(_3667__31_), .B(_3432__bF_buf4), .C(_3433__bF_buf8), .Y(_2001_) );
NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(e_reg_31_), .B(_113__bF_buf3), .Y(_2002_) );
NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf3), .B(d_reg_31_), .Y(_2003_) );
NAND3X1 NAND3X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2001_), .B(_2003_), .C(_2002_), .Y(_10__31_) );
INVX1 INVX1_880 ( .gnd(gnd), .vdd(vdd), .A(_3667__128_), .Y(_2004_) );
INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf5), .Y(_2005_) );
OAI21X1 OAI21X1_1188 ( .gnd(gnd), .vdd(vdd), .A(_3431__bF_buf2), .B(_3386__bF_buf1), .C(_2005__bF_buf11), .Y(_2006_) );
OAI21X1 OAI21X1_1189 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf10), .B(a_reg_0_), .C(_2006__bF_buf8), .Y(_2007_) );
NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(_2004_), .B(_3384_), .Y(_2008_) );
AOI22X1 AOI22X1_799 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf4), .B(_2008_), .C(_2004_), .D(_2007_), .Y(_0__0_) );
XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_3667__129_), .B(a_reg_1_), .Y(_2009_) );
XNOR2X1 XNOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(_2009_), .B(_2008_), .Y(_2010_) );
OAI22X1 OAI22X1_61 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_2006__bF_buf7), .C(_2005__bF_buf9), .D(_2010_), .Y(_0__1_) );
NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2008_), .B(_2009_), .Y(_2011_) );
OAI21X1 OAI21X1_1190 ( .gnd(gnd), .vdd(vdd), .A(_3498_), .B(_3436_), .C(_2011_), .Y(_2012_) );
NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .B(_3501_), .Y(_2013_) );
NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(_3667__130_), .B(a_reg_2_), .Y(_2014_) );
NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(_2014_), .B(_2013_), .Y(_2015_) );
XNOR2X1 XNOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2015_), .Y(_2016_) );
OAI22X1 OAI22X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3559_), .B(_2006__bF_buf6), .C(_2005__bF_buf8), .D(_2016_), .Y(_0__2_) );
AOI21X1 AOI21X1_199 ( .gnd(gnd), .vdd(vdd), .A(_2012_), .B(_2015_), .C(_2013_), .Y(_2017_) );
NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_3562_), .Y(_2018_) );
NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(_3667__131_), .B(a_reg_3_), .Y(_2019_) );
NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2019_), .B(_2018_), .Y(_2020_) );
XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(_2017_), .B(_2020_), .Y(_2021_) );
OAI22X1 OAI22X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3626_), .B(_2006__bF_buf5), .C(_2005__bF_buf7), .D(_2021_), .Y(_0__3_) );
XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_3667__132_), .B(a_reg_4_), .Y(_2022_) );
INVX1 INVX1_881 ( .gnd(gnd), .vdd(vdd), .A(_2018_), .Y(_2023_) );
OAI21X1 OAI21X1_1191 ( .gnd(gnd), .vdd(vdd), .A(_2019_), .B(_2017_), .C(_2023_), .Y(_2024_) );
XNOR2X1 XNOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(_2024_), .B(_2022_), .Y(_2025_) );
OAI22X1 OAI22X1_64 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_2006__bF_buf4), .C(_2005__bF_buf6), .D(_2025_), .Y(_0__4_) );
NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2022_), .B(_2024_), .Y(_2026_) );
OAI21X1 OAI21X1_1192 ( .gnd(gnd), .vdd(vdd), .A(_46_), .B(_3629_), .C(_2026_), .Y(_2027_) );
XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(_3667__133_), .B(a_reg_5_), .Y(_2028_) );
NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(_2027_), .Y(_2029_) );
INVX1 INVX1_882 ( .gnd(gnd), .vdd(vdd), .A(_2029_), .Y(_2030_) );
OAI21X1 OAI21X1_1193 ( .gnd(gnd), .vdd(vdd), .A(_2028_), .B(_2027_), .C(digest_valid_new_bF_buf3), .Y(_2031_) );
OAI22X1 OAI22X1_65 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_2006__bF_buf3), .C(_2031_), .D(_2030_), .Y(_0__5_) );
INVX1 INVX1_883 ( .gnd(gnd), .vdd(vdd), .A(a_reg_5_), .Y(_2032_) );
OAI21X1 OAI21X1_1194 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(_2032_), .C(_2029_), .Y(_2033_) );
AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(_3667__134_), .B(a_reg_6_), .Y(_2034_) );
NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(_3667__134_), .B(a_reg_6_), .Y(_2035_) );
NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(_2035_), .B(_2034_), .Y(_2036_) );
AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(_2033_), .B(_2036_), .Y(_2037_) );
OAI21X1 OAI21X1_1195 ( .gnd(gnd), .vdd(vdd), .A(_2036_), .B(_2033_), .C(digest_valid_new_bF_buf2), .Y(_2038_) );
OAI22X1 OAI22X1_66 ( .gnd(gnd), .vdd(vdd), .A(_181_), .B(_2006__bF_buf2), .C(_2037_), .D(_2038_), .Y(_0__6_) );
XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_3667__135_), .B(a_reg_7_), .Y(_2039_) );
OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(_2037_), .B(_2034_), .Y(_2040_) );
AOI21X1 AOI21X1_200 ( .gnd(gnd), .vdd(vdd), .A(_2040_), .B(_2039_), .C(_2005__bF_buf5), .Y(_2041_) );
OAI21X1 OAI21X1_1196 ( .gnd(gnd), .vdd(vdd), .A(_2039_), .B(_2040_), .C(_2041_), .Y(_2042_) );
OAI21X1 OAI21X1_1197 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_2006__bF_buf1), .C(_2042_), .Y(_0__7_) );
INVX1 INVX1_884 ( .gnd(gnd), .vdd(vdd), .A(a_reg_7_), .Y(_2043_) );
NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(_2034_), .B(_2039_), .Y(_2044_) );
OAI21X1 OAI21X1_1198 ( .gnd(gnd), .vdd(vdd), .A(_232_), .B(_2043_), .C(_2044_), .Y(_2045_) );
AOI21X1 AOI21X1_201 ( .gnd(gnd), .vdd(vdd), .A(_2037_), .B(_2039_), .C(_2045_), .Y(_2046_) );
INVX1 INVX1_885 ( .gnd(gnd), .vdd(vdd), .A(_3667__136_), .Y(_2047_) );
NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(_2047_), .B(_303_), .Y(_2048_) );
NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(_3667__136_), .B(a_reg_8_), .Y(_2049_) );
NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(_2049_), .B(_2048_), .Y(_2050_) );
INVX1 INVX1_886 ( .gnd(gnd), .vdd(vdd), .A(_2050_), .Y(_2051_) );
AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(_2046_), .B(_2051_), .Y(_2052_) );
OAI21X1 OAI21X1_1199 ( .gnd(gnd), .vdd(vdd), .A(_2051_), .B(_2046_), .C(digest_valid_new_bF_buf1), .Y(_2053_) );
OAI21X1 OAI21X1_1200 ( .gnd(gnd), .vdd(vdd), .A(_3667__136_), .B(_3432__bF_buf3), .C(_2005__bF_buf4), .Y(_2054_) );
OAI21X1 OAI21X1_1201 ( .gnd(gnd), .vdd(vdd), .A(_2052_), .B(_2053_), .C(_2054_), .Y(_0__8_) );
INVX1 INVX1_887 ( .gnd(gnd), .vdd(vdd), .A(_2048_), .Y(_2055_) );
OAI21X1 OAI21X1_1202 ( .gnd(gnd), .vdd(vdd), .A(_2049_), .B(_2046_), .C(_2055_), .Y(_2056_) );
XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_3667__137_), .B(a_reg_9_), .Y(_2057_) );
XNOR2X1 XNOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(_2056_), .B(_2057_), .Y(_2058_) );
OAI21X1 OAI21X1_1203 ( .gnd(gnd), .vdd(vdd), .A(_3667__137_), .B(_3432__bF_buf2), .C(_2005__bF_buf3), .Y(_2059_) );
OAI21X1 OAI21X1_1204 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf2), .B(_2058_), .C(_2059_), .Y(_0__9_) );
AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(_3667__138_), .B(a_reg_10_), .Y(_2060_) );
NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(_3667__138_), .B(a_reg_10_), .Y(_2061_) );
NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(_2061_), .B(_2060_), .Y(_2062_) );
OAI21X1 OAI21X1_1205 ( .gnd(gnd), .vdd(vdd), .A(_366_), .B(_306_), .C(_2055_), .Y(_2063_) );
OAI21X1 OAI21X1_1206 ( .gnd(gnd), .vdd(vdd), .A(_3667__137_), .B(a_reg_9_), .C(_2063_), .Y(_2064_) );
NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2057_), .B(_2050_), .Y(_2065_) );
OAI21X1 OAI21X1_1207 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_2046_), .C(_2064_), .Y(_2066_) );
AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(_2066_), .B(_2062_), .Y(_2067_) );
OAI21X1 OAI21X1_1208 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(_2066_), .C(digest_valid_new_bF_buf0), .Y(_2068_) );
OAI22X1 OAI22X1_67 ( .gnd(gnd), .vdd(vdd), .A(_438_), .B(_2006__bF_buf0), .C(_2067_), .D(_2068_), .Y(_0__10_) );
NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2060_), .B(_2067_), .Y(_2069_) );
NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_806_), .Y(_2070_) );
NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(_3667__139_), .B(a_reg_11_), .Y(_2071_) );
NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2071_), .B(_2070_), .Y(_2072_) );
XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_2069_), .B(_2072_), .Y(_2073_) );
OAI22X1 OAI22X1_68 ( .gnd(gnd), .vdd(vdd), .A(_503_), .B(_2006__bF_buf8), .C(_2005__bF_buf1), .D(_2073_), .Y(_0__11_) );
NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_2062_), .B(_2072_), .Y(_2074_) );
NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2065_), .B(_2074_), .Y(_2075_) );
INVX1 INVX1_888 ( .gnd(gnd), .vdd(vdd), .A(_2075_), .Y(_2076_) );
AOI21X1 AOI21X1_202 ( .gnd(gnd), .vdd(vdd), .A(_2072_), .B(_2060_), .C(_2070_), .Y(_2077_) );
OAI21X1 OAI21X1_1209 ( .gnd(gnd), .vdd(vdd), .A(_2074_), .B(_2064_), .C(_2077_), .Y(_2078_) );
INVX1 INVX1_889 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .Y(_2079_) );
OAI21X1 OAI21X1_1210 ( .gnd(gnd), .vdd(vdd), .A(_2076_), .B(_2046_), .C(_2079_), .Y(_2080_) );
AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(_3667__140_), .B(a_reg_12_), .Y(_2081_) );
NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(_3667__140_), .B(a_reg_12_), .Y(_2082_) );
NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2082_), .B(_2081_), .Y(_2083_) );
AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(_2080_), .B(_2083_), .Y(_2084_) );
OAI21X1 OAI21X1_1211 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_2080_), .C(digest_valid_new_bF_buf8), .Y(_2085_) );
OAI22X1 OAI22X1_69 ( .gnd(gnd), .vdd(vdd), .A(_570_), .B(_2006__bF_buf7), .C(_2084_), .D(_2085_), .Y(_0__12_) );
NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2081_), .B(_2084_), .Y(_2086_) );
NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(_635_), .B(_918_), .Y(_2087_) );
NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(_3667__141_), .B(a_reg_13_), .Y(_2088_) );
NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .B(_2087_), .Y(_2089_) );
XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(_2086_), .B(_2089_), .Y(_2090_) );
OAI21X1 OAI21X1_1212 ( .gnd(gnd), .vdd(vdd), .A(_3667__141_), .B(_3432__bF_buf1), .C(_2005__bF_buf0), .Y(_2091_) );
OAI21X1 OAI21X1_1213 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf11), .B(_2090_), .C(_2091_), .Y(_0__13_) );
INVX1 INVX1_890 ( .gnd(gnd), .vdd(vdd), .A(a_reg_14_), .Y(_2092_) );
NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_2092_), .Y(_2093_) );
NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(_3667__142_), .B(a_reg_14_), .Y(_2094_) );
NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(_2094_), .B(_2093_), .Y(_2095_) );
INVX1 INVX1_891 ( .gnd(gnd), .vdd(vdd), .A(_2095_), .Y(_2096_) );
INVX1 INVX1_892 ( .gnd(gnd), .vdd(vdd), .A(_2088_), .Y(_2097_) );
OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(_2087_), .B(_2081_), .Y(_2098_) );
OAI21X1 OAI21X1_1214 ( .gnd(gnd), .vdd(vdd), .A(_2098_), .B(_2084_), .C(_2097_), .Y(_2099_) );
OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(_2099_), .B(_2096_), .Y(_2100_) );
OAI21X1 OAI21X1_1215 ( .gnd(gnd), .vdd(vdd), .A(_2093_), .B(_2094_), .C(_2099_), .Y(_2101_) );
NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_2101_), .B(_2100_), .Y(_2102_) );
OAI22X1 OAI22X1_70 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_2006__bF_buf6), .C(_2005__bF_buf10), .D(_2102_), .Y(_0__14_) );
OAI21X1 OAI21X1_1216 ( .gnd(gnd), .vdd(vdd), .A(_699_), .B(_2092_), .C(_2100_), .Y(_2103_) );
AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(_3667__143_), .B(a_reg_15_), .Y(_2104_) );
NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3667__143_), .B(a_reg_15_), .Y(_2105_) );
NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(_2105_), .B(_2104_), .Y(_2106_) );
XNOR2X1 XNOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(_2103_), .B(_2106_), .Y(_2107_) );
OAI22X1 OAI22X1_71 ( .gnd(gnd), .vdd(vdd), .A(_769_), .B(_2006__bF_buf5), .C(_2005__bF_buf9), .D(_2107_), .Y(_0__15_) );
OAI21X1 OAI21X1_1217 ( .gnd(gnd), .vdd(vdd), .A(_3667__141_), .B(a_reg_13_), .C(_2098_), .Y(_2108_) );
AOI21X1 AOI21X1_203 ( .gnd(gnd), .vdd(vdd), .A(_2106_), .B(_2093_), .C(_2104_), .Y(_2109_) );
NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_2106_), .B(_2095_), .Y(_2110_) );
OAI21X1 OAI21X1_1218 ( .gnd(gnd), .vdd(vdd), .A(_2110_), .B(_2108_), .C(_2109_), .Y(_2111_) );
NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(_2083_), .B(_2089_), .Y(_2112_) );
NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(_2112_), .B(_2110_), .Y(_2113_) );
AOI21X1 AOI21X1_204 ( .gnd(gnd), .vdd(vdd), .A(_2078_), .B(_2113_), .C(_2111_), .Y(_2114_) );
NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2075_), .B(_2113_), .Y(_2115_) );
OAI21X1 OAI21X1_1219 ( .gnd(gnd), .vdd(vdd), .A(_2115_), .B(_2046_), .C(_2114_), .Y(_2116_) );
INVX1 INVX1_893 ( .gnd(gnd), .vdd(vdd), .A(a_reg_16_), .Y(_2117_) );
NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_2117_), .Y(_2118_) );
NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(_3667__144_), .B(a_reg_16_), .Y(_2119_) );
NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(_2119_), .B(_2118_), .Y(_2120_) );
NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_2116_), .Y(_2121_) );
NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_2116_), .Y(_2122_) );
NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf7), .B(_2122_), .Y(_2123_) );
OAI21X1 OAI21X1_1220 ( .gnd(gnd), .vdd(vdd), .A(_3667__144_), .B(_3432__bF_buf0), .C(_2005__bF_buf8), .Y(_2124_) );
OAI21X1 OAI21X1_1221 ( .gnd(gnd), .vdd(vdd), .A(_2121_), .B(_2123_), .C(_2124_), .Y(_0__16_) );
NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_843_), .Y(_2125_) );
NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(_3667__145_), .B(a_reg_17_), .Y(_2126_) );
NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(_2126_), .B(_2125_), .Y(_2127_) );
OAI21X1 OAI21X1_1222 ( .gnd(gnd), .vdd(vdd), .A(_840_), .B(_2117_), .C(_2122_), .Y(_2128_) );
XNOR2X1 XNOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(_2128_), .B(_2127_), .Y(_2129_) );
OAI22X1 OAI22X1_72 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_2006__bF_buf4), .C(_2005__bF_buf7), .D(_2129_), .Y(_0__17_) );
AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(_2120_), .B(_2127_), .Y(_2130_) );
NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(_2118_), .B(_2127_), .Y(_2131_) );
OAI21X1 OAI21X1_1223 ( .gnd(gnd), .vdd(vdd), .A(_894_), .B(_843_), .C(_2131_), .Y(_2132_) );
AOI21X1 AOI21X1_205 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2130_), .C(_2132_), .Y(_2133_) );
NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1214_), .Y(_2134_) );
NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(_3667__146_), .B(a_reg_18_), .Y(_2135_) );
OAI21X1 OAI21X1_1224 ( .gnd(gnd), .vdd(vdd), .A(_2134_), .B(_2135_), .C(_2133_), .Y(_2136_) );
NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(_2135_), .B(_2134_), .Y(_2137_) );
INVX1 INVX1_894 ( .gnd(gnd), .vdd(vdd), .A(_2137_), .Y(_2138_) );
OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(_2133_), .B(_2138_), .Y(_2139_) );
NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2136_), .B(_2139_), .Y(_2140_) );
OAI21X1 OAI21X1_1225 ( .gnd(gnd), .vdd(vdd), .A(_3667__146_), .B(_3432__bF_buf11), .C(_2005__bF_buf6), .Y(_2141_) );
OAI21X1 OAI21X1_1226 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf5), .B(_2140_), .C(_2141_), .Y(_0__18_) );
OAI21X1 OAI21X1_1227 ( .gnd(gnd), .vdd(vdd), .A(_941_), .B(_1214_), .C(_2139_), .Y(_2142_) );
XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_3667__147_), .B(a_reg_19_), .Y(_2143_) );
OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(_2142_), .B(_2143_), .Y(_2144_) );
NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2142_), .Y(_2145_) );
NAND3X1 NAND3X1_294 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf6), .B(_2145_), .C(_2144_), .Y(_2146_) );
OAI21X1 OAI21X1_1228 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .B(_2006__bF_buf3), .C(_2146_), .Y(_0__19_) );
NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_2143_), .B(_2137_), .Y(_2147_) );
INVX1 INVX1_895 ( .gnd(gnd), .vdd(vdd), .A(_2147_), .Y(_2148_) );
NAND3X1 NAND3X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2130_), .B(_2148_), .C(_2116_), .Y(_2149_) );
OAI21X1 OAI21X1_1229 ( .gnd(gnd), .vdd(vdd), .A(_3667__147_), .B(a_reg_19_), .C(_2134_), .Y(_2150_) );
OAI21X1 OAI21X1_1230 ( .gnd(gnd), .vdd(vdd), .A(_1003_), .B(_1279_), .C(_2150_), .Y(_2151_) );
AOI21X1 AOI21X1_206 ( .gnd(gnd), .vdd(vdd), .A(_2132_), .B(_2148_), .C(_2151_), .Y(_2152_) );
AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(_2149_), .B(_2152_), .Y(_2153_) );
NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_1358_), .Y(_2154_) );
NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(_3667__148_), .B(a_reg_20_), .Y(_2155_) );
NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(_2155_), .B(_2154_), .Y(_2156_) );
INVX1 INVX1_896 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .Y(_2157_) );
NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(_2157_), .B(_2153_), .Y(_2158_) );
INVX1 INVX1_897 ( .gnd(gnd), .vdd(vdd), .A(_2153_), .Y(_2159_) );
OAI21X1 OAI21X1_1231 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .B(_2159_), .C(digest_valid_new_bF_buf5), .Y(_2160_) );
OAI22X1 OAI22X1_73 ( .gnd(gnd), .vdd(vdd), .A(_1072_), .B(_2006__bF_buf2), .C(_2158_), .D(_2160_), .Y(_0__20_) );
NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_1362_), .Y(_2161_) );
NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(_3667__149_), .B(a_reg_21_), .Y(_2162_) );
NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(_2162_), .B(_2161_), .Y(_2163_) );
NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(_2154_), .B(_2158_), .Y(_2164_) );
XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(_2164_), .B(_2163_), .Y(_2165_) );
OAI22X1 OAI22X1_74 ( .gnd(gnd), .vdd(vdd), .A(_1128_), .B(_2006__bF_buf1), .C(_2005__bF_buf4), .D(_2165_), .Y(_0__21_) );
NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .B(_2163_), .Y(_2166_) );
AOI21X1 AOI21X1_207 ( .gnd(gnd), .vdd(vdd), .A(_2163_), .B(_2154_), .C(_2161_), .Y(_2167_) );
OAI21X1 OAI21X1_1232 ( .gnd(gnd), .vdd(vdd), .A(_2166_), .B(_2153_), .C(_2167_), .Y(_2168_) );
NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1405_), .Y(_2169_) );
NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(_3667__150_), .B(a_reg_22_), .Y(_2170_) );
NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(_2170_), .B(_2169_), .Y(_2171_) );
NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2168_), .Y(_2172_) );
NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2168_), .Y(_2173_) );
NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf4), .B(_2173_), .Y(_2174_) );
OAI21X1 OAI21X1_1233 ( .gnd(gnd), .vdd(vdd), .A(_3667__150_), .B(_3432__bF_buf10), .C(_2005__bF_buf3), .Y(_2175_) );
OAI21X1 OAI21X1_1234 ( .gnd(gnd), .vdd(vdd), .A(_2172_), .B(_2174_), .C(_2175_), .Y(_0__22_) );
OAI21X1 OAI21X1_1235 ( .gnd(gnd), .vdd(vdd), .A(_1188_), .B(_1405_), .C(_2173_), .Y(_2176_) );
XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_3667__151_), .B(a_reg_23_), .Y(_2177_) );
NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_2177_), .B(_2176_), .Y(_2178_) );
OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(_2176_), .B(_2177_), .Y(_2179_) );
NAND3X1 NAND3X1_296 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf3), .B(_2178_), .C(_2179_), .Y(_2180_) );
OAI21X1 OAI21X1_1236 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_2006__bF_buf0), .C(_2180_), .Y(_0__23_) );
INVX1 INVX1_898 ( .gnd(gnd), .vdd(vdd), .A(_2167_), .Y(_2181_) );
AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(_2171_), .B(_2177_), .Y(_2182_) );
OAI21X1 OAI21X1_1237 ( .gnd(gnd), .vdd(vdd), .A(_3667__151_), .B(a_reg_23_), .C(_2169_), .Y(_2183_) );
OAI21X1 OAI21X1_1238 ( .gnd(gnd), .vdd(vdd), .A(_1244_), .B(_1483_), .C(_2183_), .Y(_2184_) );
AOI21X1 AOI21X1_208 ( .gnd(gnd), .vdd(vdd), .A(_2181_), .B(_2182_), .C(_2184_), .Y(_2185_) );
NAND3X1 NAND3X1_297 ( .gnd(gnd), .vdd(vdd), .A(_2156_), .B(_2163_), .C(_2182_), .Y(_2186_) );
OAI21X1 OAI21X1_1239 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2152_), .C(_2185_), .Y(_2187_) );
NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(_2130_), .B(_2148_), .Y(_2188_) );
NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(_2186_), .B(_2188_), .Y(_2189_) );
AOI21X1 AOI21X1_209 ( .gnd(gnd), .vdd(vdd), .A(_2116_), .B(_2189_), .C(_2187_), .Y(_2190_) );
INVX1 INVX1_899 ( .gnd(gnd), .vdd(vdd), .A(_3667__152_), .Y(_2191_) );
NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(_2191_), .B(_1247_), .Y(_2192_) );
NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(_3667__152_), .B(a_reg_24_), .Y(_2193_) );
NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2192_), .Y(_2194_) );
INVX1 INVX1_900 ( .gnd(gnd), .vdd(vdd), .A(_2194_), .Y(_2195_) );
AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(_2190_), .B(_2195_), .Y(_2196_) );
OAI21X1 OAI21X1_1240 ( .gnd(gnd), .vdd(vdd), .A(_2195_), .B(_2190_), .C(digest_valid_new_bF_buf2), .Y(_2197_) );
OAI21X1 OAI21X1_1241 ( .gnd(gnd), .vdd(vdd), .A(_3667__152_), .B(_3432__bF_buf9), .C(_2005__bF_buf2), .Y(_2198_) );
OAI21X1 OAI21X1_1242 ( .gnd(gnd), .vdd(vdd), .A(_2196_), .B(_2197_), .C(_2198_), .Y(_0__24_) );
INVX1 INVX1_901 ( .gnd(gnd), .vdd(vdd), .A(_2192_), .Y(_2199_) );
OAI21X1 OAI21X1_1243 ( .gnd(gnd), .vdd(vdd), .A(_2193_), .B(_2190_), .C(_2199_), .Y(_2200_) );
NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(_1331_), .B(_1538_), .Y(_2201_) );
NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(_3667__153_), .B(a_reg_25_), .Y(_2202_) );
NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(_2202_), .B(_2201_), .Y(_2203_) );
XNOR2X1 XNOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(_2200_), .B(_2203_), .Y(_2204_) );
OAI21X1 OAI21X1_1244 ( .gnd(gnd), .vdd(vdd), .A(_3667__153_), .B(_3432__bF_buf8), .C(_2005__bF_buf1), .Y(_2205_) );
OAI21X1 OAI21X1_1245 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf0), .B(_2204_), .C(_2205_), .Y(_0__25_) );
INVX1 INVX1_902 ( .gnd(gnd), .vdd(vdd), .A(_2203_), .Y(_2206_) );
NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2195_), .B(_2206_), .Y(_2207_) );
INVX1 INVX1_903 ( .gnd(gnd), .vdd(vdd), .A(_2207_), .Y(_2208_) );
AOI21X1 AOI21X1_210 ( .gnd(gnd), .vdd(vdd), .A(_2203_), .B(_2192_), .C(_2201_), .Y(_2209_) );
OAI21X1 OAI21X1_1246 ( .gnd(gnd), .vdd(vdd), .A(_2208_), .B(_2190_), .C(_2209_), .Y(_2210_) );
INVX1 INVX1_904 ( .gnd(gnd), .vdd(vdd), .A(a_reg_26_), .Y(_2211_) );
NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .B(_2211_), .Y(_2212_) );
NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(_3667__154_), .B(a_reg_26_), .Y(_2213_) );
NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2213_), .B(_2212_), .Y(_2214_) );
NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2210_), .Y(_2215_) );
NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2210_), .Y(_2216_) );
NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf1), .B(_2216_), .Y(_2217_) );
OAI21X1 OAI21X1_1247 ( .gnd(gnd), .vdd(vdd), .A(_3667__154_), .B(_3432__bF_buf7), .C(_2005__bF_buf11), .Y(_2218_) );
OAI21X1 OAI21X1_1248 ( .gnd(gnd), .vdd(vdd), .A(_2215_), .B(_2217_), .C(_2218_), .Y(_0__26_) );
XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(a_reg_27_), .B(_3667__155_), .Y(_2219_) );
OAI21X1 OAI21X1_1249 ( .gnd(gnd), .vdd(vdd), .A(_1381_), .B(_2211_), .C(_2216_), .Y(_2220_) );
XNOR2X1 XNOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(_2220_), .B(_2219_), .Y(_2221_) );
OAI22X1 OAI22X1_75 ( .gnd(gnd), .vdd(vdd), .A(_1422_), .B(_2006__bF_buf8), .C(_2005__bF_buf10), .D(_2221_), .Y(_0__27_) );
INVX1 INVX1_905 ( .gnd(gnd), .vdd(vdd), .A(_2209_), .Y(_2222_) );
AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(_2214_), .B(_2219_), .Y(_2223_) );
INVX1 INVX1_906 ( .gnd(gnd), .vdd(vdd), .A(a_reg_27_), .Y(_2224_) );
NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_2212_), .B(_2219_), .Y(_2225_) );
OAI21X1 OAI21X1_1250 ( .gnd(gnd), .vdd(vdd), .A(_2224_), .B(_1422_), .C(_2225_), .Y(_2226_) );
AOI21X1 AOI21X1_211 ( .gnd(gnd), .vdd(vdd), .A(_2222_), .B(_2223_), .C(_2226_), .Y(_2227_) );
NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(_2223_), .B(_2207_), .Y(_2228_) );
OAI21X1 OAI21X1_1251 ( .gnd(gnd), .vdd(vdd), .A(_2228_), .B(_2190_), .C(_2227_), .Y(_2229_) );
NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(a_reg_28_), .B(_3667__156_), .Y(_2230_) );
OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(a_reg_28_), .B(_3667__156_), .Y(_2231_) );
NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_2230_), .B(_2231_), .Y(_2232_) );
XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_2232_), .Y(_2233_) );
OAI22X1 OAI22X1_76 ( .gnd(gnd), .vdd(vdd), .A(_1467_), .B(_2006__bF_buf7), .C(_2005__bF_buf9), .D(_2233_), .Y(_0__28_) );
INVX1 INVX1_907 ( .gnd(gnd), .vdd(vdd), .A(_1503_), .Y(_2234_) );
INVX1 INVX1_908 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .Y(_2235_) );
OAI21X1 OAI21X1_1252 ( .gnd(gnd), .vdd(vdd), .A(_2232_), .B(_2235_), .C(_2230_), .Y(_2236_) );
INVX1 INVX1_909 ( .gnd(gnd), .vdd(vdd), .A(a_reg_29_), .Y(_2237_) );
NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2237_), .B(_1502_), .Y(_2238_) );
NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(a_reg_29_), .B(_3667__157_), .Y(_2239_) );
NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(_2239_), .B(_2238_), .Y(_2240_) );
INVX1 INVX1_910 ( .gnd(gnd), .vdd(vdd), .A(_2240_), .Y(_2241_) );
OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(_2236_), .B(_2241_), .Y(_2242_) );
AOI21X1 AOI21X1_212 ( .gnd(gnd), .vdd(vdd), .A(_2236_), .B(_2241_), .C(_2005__bF_buf8), .Y(_2243_) );
AOI22X1 AOI22X1_800 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf7), .B(_2234_), .C(_2243_), .D(_2242_), .Y(_0__29_) );
XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(a_reg_30_), .B(_3667__158_), .Y(_2244_) );
INVX1 INVX1_911 ( .gnd(gnd), .vdd(vdd), .A(_2244_), .Y(_2245_) );
INVX1 INVX1_912 ( .gnd(gnd), .vdd(vdd), .A(_2238_), .Y(_2246_) );
OAI21X1 OAI21X1_1253 ( .gnd(gnd), .vdd(vdd), .A(_2230_), .B(_2239_), .C(_2246_), .Y(_2247_) );
NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(_2232_), .B(_2241_), .Y(_2248_) );
AOI21X1 AOI21X1_213 ( .gnd(gnd), .vdd(vdd), .A(_2229_), .B(_2248_), .C(_2247_), .Y(_2249_) );
AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(_2249_), .B(_2245_), .Y(_2250_) );
OAI21X1 OAI21X1_1254 ( .gnd(gnd), .vdd(vdd), .A(_2245_), .B(_2249_), .C(digest_valid_new_bF_buf0), .Y(_2251_) );
OAI21X1 OAI21X1_1255 ( .gnd(gnd), .vdd(vdd), .A(_3667__158_), .B(_3432__bF_buf6), .C(_2005__bF_buf6), .Y(_2252_) );
OAI21X1 OAI21X1_1256 ( .gnd(gnd), .vdd(vdd), .A(_2250_), .B(_2251_), .C(_2252_), .Y(_0__30_) );
NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(a_reg_30_), .B(_3667__158_), .Y(_2253_) );
OAI21X1 OAI21X1_1257 ( .gnd(gnd), .vdd(vdd), .A(_2245_), .B(_2249_), .C(_2253_), .Y(_2254_) );
XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(a_reg_31_), .B(_3667__159_), .Y(_2255_) );
NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_2255_), .B(_2254_), .Y(_2256_) );
OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(_2254_), .B(_2255_), .Y(_2257_) );
NAND3X1 NAND3X1_298 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(_2256_), .C(_2257_), .Y(_2258_) );
OAI21X1 OAI21X1_1258 ( .gnd(gnd), .vdd(vdd), .A(_1592_), .B(_2006__bF_buf6), .C(_2258_), .Y(_0__31_) );
NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(b_reg_0_), .B(_3667__96_), .Y(_2259_) );
OAI21X1 OAI21X1_1259 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_1595_), .C(digest_valid_new_bF_buf7), .Y(_2260_) );
OAI21X1 OAI21X1_1260 ( .gnd(gnd), .vdd(vdd), .A(_3667__96_), .B(_3432__bF_buf5), .C(_2005__bF_buf5), .Y(_2261_) );
OAI21X1 OAI21X1_1261 ( .gnd(gnd), .vdd(vdd), .A(_2259_), .B(_2260_), .C(_2261_), .Y(_1__0_) );
NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(_3412_), .B(_1595_), .Y(_2262_) );
XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(b_reg_1_), .B(_3667__97_), .Y(_2263_) );
XNOR2X1 XNOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(_2263_), .B(_2262_), .Y(_2264_) );
OAI22X1 OAI22X1_77 ( .gnd(gnd), .vdd(vdd), .A(_1598_), .B(_2006__bF_buf5), .C(_2005__bF_buf4), .D(_2264_), .Y(_1__1_) );
NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2262_), .B(_2263_), .Y(_2265_) );
OAI21X1 OAI21X1_1262 ( .gnd(gnd), .vdd(vdd), .A(_3440_), .B(_1598_), .C(_2265_), .Y(_2266_) );
NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(_1601_), .B(_1602_), .Y(_2267_) );
NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(b_reg_2_), .B(_3667__98_), .Y(_2268_) );
NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(_2268_), .B(_2267_), .Y(_2269_) );
XNOR2X1 XNOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(_2266_), .B(_2269_), .Y(_2270_) );
OAI22X1 OAI22X1_78 ( .gnd(gnd), .vdd(vdd), .A(_1602_), .B(_2006__bF_buf4), .C(_2005__bF_buf3), .D(_2270_), .Y(_1__2_) );
AOI21X1 AOI21X1_214 ( .gnd(gnd), .vdd(vdd), .A(_2266_), .B(_2269_), .C(_2267_), .Y(_2271_) );
NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(_3575_), .B(_1605_), .Y(_2272_) );
NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(b_reg_3_), .B(_3667__99_), .Y(_2273_) );
NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(_2273_), .B(_2272_), .Y(_2274_) );
XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_2271_), .B(_2274_), .Y(_2275_) );
OAI21X1 OAI21X1_1263 ( .gnd(gnd), .vdd(vdd), .A(_3667__99_), .B(_3432__bF_buf4), .C(_2005__bF_buf2), .Y(_2276_) );
OAI21X1 OAI21X1_1264 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf1), .B(_2275_), .C(_2276_), .Y(_1__3_) );
NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(b_reg_4_), .B(_3667__100_), .Y(_2277_) );
NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_3642_), .B(_1608_), .Y(_2278_) );
NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(_2277_), .B(_2278_), .Y(_2279_) );
OAI21X1 OAI21X1_1265 ( .gnd(gnd), .vdd(vdd), .A(_3575_), .B(_1605_), .C(_2271_), .Y(_2280_) );
OAI21X1 OAI21X1_1266 ( .gnd(gnd), .vdd(vdd), .A(b_reg_3_), .B(_3667__99_), .C(_2280_), .Y(_2281_) );
XNOR2X1 XNOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(_2281_), .B(_2279_), .Y(_2282_) );
OAI22X1 OAI22X1_79 ( .gnd(gnd), .vdd(vdd), .A(_1608_), .B(_2006__bF_buf3), .C(_2005__bF_buf0), .D(_2282_), .Y(_1__4_) );
OAI21X1 OAI21X1_1267 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2281_), .C(_2277_), .Y(_2283_) );
NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(b_reg_5_), .B(_3667__101_), .Y(_2284_) );
INVX1 INVX1_913 ( .gnd(gnd), .vdd(vdd), .A(_2284_), .Y(_2285_) );
NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(b_reg_5_), .B(_3667__101_), .Y(_2286_) );
OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(_2285_), .B(_2286_), .Y(_2287_) );
INVX1 INVX1_914 ( .gnd(gnd), .vdd(vdd), .A(_2287_), .Y(_2288_) );
NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2288_), .B(_2283_), .Y(_2289_) );
INVX1 INVX1_915 ( .gnd(gnd), .vdd(vdd), .A(_2289_), .Y(_2290_) );
OAI21X1 OAI21X1_1268 ( .gnd(gnd), .vdd(vdd), .A(_2288_), .B(_2283_), .C(digest_valid_new_bF_buf6), .Y(_2291_) );
OAI22X1 OAI22X1_80 ( .gnd(gnd), .vdd(vdd), .A(_1611_), .B(_2006__bF_buf2), .C(_2291_), .D(_2290_), .Y(_1__5_) );
OAI21X1 OAI21X1_1269 ( .gnd(gnd), .vdd(vdd), .A(_60_), .B(_1611_), .C(_2289_), .Y(_2292_) );
NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .B(_1615_), .Y(_2293_) );
INVX1 INVX1_916 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .Y(_2294_) );
NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_1614_), .B(_1615_), .Y(_2295_) );
NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(_2295_), .B(_2294_), .Y(_2296_) );
XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(_2292_), .B(_2296_), .Y(_2297_) );
OAI22X1 OAI22X1_81 ( .gnd(gnd), .vdd(vdd), .A(_1615_), .B(_2006__bF_buf1), .C(_2005__bF_buf11), .D(_2297_), .Y(_1__6_) );
AOI21X1 AOI21X1_215 ( .gnd(gnd), .vdd(vdd), .A(_2292_), .B(_2295_), .C(_2293_), .Y(_2298_) );
NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(b_reg_7_), .B(_3667__103_), .Y(_2299_) );
NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(b_reg_7_), .B(_3667__103_), .Y(_2300_) );
INVX1 INVX1_917 ( .gnd(gnd), .vdd(vdd), .A(_2300_), .Y(_2301_) );
NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .B(_2301_), .Y(_2302_) );
INVX1 INVX1_918 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .Y(_2303_) );
NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(_2303_), .B(_2298_), .Y(_2304_) );
INVX1 INVX1_919 ( .gnd(gnd), .vdd(vdd), .A(_2304_), .Y(_2305_) );
NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(_2303_), .B(_2298_), .Y(_2306_) );
OAI21X1 OAI21X1_1270 ( .gnd(gnd), .vdd(vdd), .A(_2306_), .B(_2305_), .C(digest_valid_new_bF_buf5), .Y(_2307_) );
OAI21X1 OAI21X1_1271 ( .gnd(gnd), .vdd(vdd), .A(_3667__103_), .B(_3432__bF_buf3), .C(_2005__bF_buf10), .Y(_2308_) );
NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_2308_), .B(_2307_), .Y(_1__7_) );
NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(_1620_), .B(_1621_), .Y(_2309_) );
NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(b_reg_8_), .B(_3667__104_), .Y(_2310_) );
NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2293_), .B(_2303_), .Y(_2311_) );
OAI21X1 OAI21X1_1272 ( .gnd(gnd), .vdd(vdd), .A(_2277_), .B(_2286_), .C(_2284_), .Y(_2312_) );
NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(_2302_), .B(_2296_), .Y(_2313_) );
NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_2312_), .B(_2313_), .Y(_2314_) );
NAND3X1 NAND3X1_299 ( .gnd(gnd), .vdd(vdd), .A(_2299_), .B(_2311_), .C(_2314_), .Y(_2315_) );
NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(_2279_), .B(_2287_), .Y(_2316_) );
NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(_2316_), .B(_2313_), .Y(_2317_) );
NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(_2317_), .B(_2281_), .Y(_2318_) );
NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(_2315_), .B(_2318_), .Y(_2319_) );
OAI21X1 OAI21X1_1273 ( .gnd(gnd), .vdd(vdd), .A(_2309_), .B(_2310_), .C(_2319_), .Y(_2320_) );
NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(_2310_), .B(_2309_), .Y(_2321_) );
OAI21X1 OAI21X1_1274 ( .gnd(gnd), .vdd(vdd), .A(_2315_), .B(_2318_), .C(_2321_), .Y(_2322_) );
NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2322_), .B(_2320_), .Y(_2323_) );
OAI21X1 OAI21X1_1275 ( .gnd(gnd), .vdd(vdd), .A(_3667__104_), .B(_3432__bF_buf2), .C(_2005__bF_buf9), .Y(_2324_) );
OAI21X1 OAI21X1_1276 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf8), .B(_2323_), .C(_2324_), .Y(_1__8_) );
OAI21X1 OAI21X1_1277 ( .gnd(gnd), .vdd(vdd), .A(_1620_), .B(_1621_), .C(_2322_), .Y(_2325_) );
XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(b_reg_9_), .B(_3667__105_), .Y(_2326_) );
XNOR2X1 XNOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(_2325_), .B(_2326_), .Y(_2327_) );
OAI21X1 OAI21X1_1278 ( .gnd(gnd), .vdd(vdd), .A(_3667__105_), .B(_3432__bF_buf1), .C(_2005__bF_buf7), .Y(_2328_) );
OAI21X1 OAI21X1_1279 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf6), .B(_2327_), .C(_2328_), .Y(_1__9_) );
NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(_1627_), .B(_1628_), .Y(_2329_) );
NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(b_reg_10_), .B(_3667__106_), .Y(_2330_) );
NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(_2330_), .B(_2329_), .Y(_2331_) );
NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_1624_), .Y(_2332_) );
AOI21X1 AOI21X1_216 ( .gnd(gnd), .vdd(vdd), .A(_2326_), .B(_2309_), .C(_2332_), .Y(_2333_) );
NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2326_), .B(_2321_), .Y(_2334_) );
OAI21X1 OAI21X1_1280 ( .gnd(gnd), .vdd(vdd), .A(_2334_), .B(_2319_), .C(_2333_), .Y(_2335_) );
AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(_2335_), .B(_2331_), .Y(_2336_) );
OAI21X1 OAI21X1_1281 ( .gnd(gnd), .vdd(vdd), .A(_2331_), .B(_2335_), .C(digest_valid_new_bF_buf4), .Y(_2337_) );
OAI22X1 OAI22X1_82 ( .gnd(gnd), .vdd(vdd), .A(_1628_), .B(_2006__bF_buf0), .C(_2336_), .D(_2337_), .Y(_1__10_) );
NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(_2329_), .B(_2336_), .Y(_2338_) );
NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(_1631_), .B(_1632_), .Y(_2339_) );
NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(b_reg_11_), .B(_3667__107_), .Y(_2340_) );
NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(_2340_), .B(_2339_), .Y(_2341_) );
XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(_2338_), .B(_2341_), .Y(_2342_) );
OAI21X1 OAI21X1_1282 ( .gnd(gnd), .vdd(vdd), .A(_3667__107_), .B(_3432__bF_buf0), .C(_2005__bF_buf5), .Y(_2343_) );
OAI21X1 OAI21X1_1283 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf4), .B(_2342_), .C(_2343_), .Y(_1__11_) );
NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2331_), .B(_2341_), .Y(_2344_) );
NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(_2334_), .B(_2344_), .Y(_2345_) );
OAI21X1 OAI21X1_1284 ( .gnd(gnd), .vdd(vdd), .A(_2315_), .B(_2318_), .C(_2345_), .Y(_2346_) );
AOI21X1 AOI21X1_217 ( .gnd(gnd), .vdd(vdd), .A(_2341_), .B(_2329_), .C(_2339_), .Y(_2347_) );
OAI21X1 OAI21X1_1285 ( .gnd(gnd), .vdd(vdd), .A(_2344_), .B(_2333_), .C(_2347_), .Y(_2348_) );
INVX1 INVX1_920 ( .gnd(gnd), .vdd(vdd), .A(_2348_), .Y(_2349_) );
AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(_2346_), .B(_2349_), .Y(_2350_) );
INVX1 INVX1_921 ( .gnd(gnd), .vdd(vdd), .A(_2350_), .Y(_2351_) );
NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(_1635_), .B(_1636_), .Y(_2352_) );
NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(b_reg_12_), .B(_3667__108_), .Y(_2353_) );
NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(_2353_), .B(_2352_), .Y(_2354_) );
AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(_2351_), .B(_2354_), .Y(_2355_) );
OAI21X1 OAI21X1_1286 ( .gnd(gnd), .vdd(vdd), .A(_2354_), .B(_2351_), .C(digest_valid_new_bF_buf3), .Y(_2356_) );
OAI22X1 OAI22X1_83 ( .gnd(gnd), .vdd(vdd), .A(_1636_), .B(_2006__bF_buf8), .C(_2355_), .D(_2356_), .Y(_1__12_) );
INVX1 INVX1_922 ( .gnd(gnd), .vdd(vdd), .A(_2352_), .Y(_2357_) );
OAI21X1 OAI21X1_1287 ( .gnd(gnd), .vdd(vdd), .A(_2353_), .B(_2350_), .C(_2357_), .Y(_2358_) );
INVX1 INVX1_923 ( .gnd(gnd), .vdd(vdd), .A(_2358_), .Y(_2359_) );
NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(_1639_), .B(_1640_), .Y(_2360_) );
NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(b_reg_13_), .B(_3667__109_), .Y(_2361_) );
NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(_2361_), .B(_2360_), .Y(_2362_) );
AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(_2359_), .B(_2362_), .Y(_2363_) );
NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(_2362_), .B(_2359_), .Y(_2364_) );
OAI21X1 OAI21X1_1288 ( .gnd(gnd), .vdd(vdd), .A(_2364_), .B(_2363_), .C(digest_valid_new_bF_buf2), .Y(_2365_) );
OAI21X1 OAI21X1_1289 ( .gnd(gnd), .vdd(vdd), .A(_3667__109_), .B(_3432__bF_buf11), .C(_2005__bF_buf3), .Y(_2366_) );
NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_2366_), .B(_2365_), .Y(_1__13_) );
AOI21X1 AOI21X1_218 ( .gnd(gnd), .vdd(vdd), .A(_2362_), .B(_2352_), .C(_2360_), .Y(_2367_) );
NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(_2354_), .B(_2362_), .Y(_2368_) );
OAI21X1 OAI21X1_1290 ( .gnd(gnd), .vdd(vdd), .A(_2368_), .B(_2350_), .C(_2367_), .Y(_2369_) );
NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1644_), .Y(_2370_) );
NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(b_reg_14_), .B(_3667__110_), .Y(_2371_) );
NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(_2371_), .B(_2370_), .Y(_2372_) );
NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2369_), .Y(_2373_) );
INVX1 INVX1_924 ( .gnd(gnd), .vdd(vdd), .A(_2373_), .Y(_2374_) );
OAI21X1 OAI21X1_1291 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2369_), .C(digest_valid_new_bF_buf1), .Y(_2375_) );
OAI22X1 OAI22X1_84 ( .gnd(gnd), .vdd(vdd), .A(_1644_), .B(_2006__bF_buf7), .C(_2375_), .D(_2374_), .Y(_1__14_) );
OAI21X1 OAI21X1_1292 ( .gnd(gnd), .vdd(vdd), .A(_1643_), .B(_1644_), .C(_2373_), .Y(_2376_) );
NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(_709_), .B(_1647_), .Y(_2377_) );
NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(b_reg_15_), .B(_3667__111_), .Y(_2378_) );
NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(_2378_), .B(_2377_), .Y(_2379_) );
XNOR2X1 XNOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(_2376_), .B(_2379_), .Y(_2380_) );
OAI21X1 OAI21X1_1293 ( .gnd(gnd), .vdd(vdd), .A(_3667__111_), .B(_3432__bF_buf10), .C(_2005__bF_buf2), .Y(_2381_) );
OAI21X1 OAI21X1_1294 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf1), .B(_2380_), .C(_2381_), .Y(_1__15_) );
NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_2372_), .B(_2379_), .Y(_2382_) );
AOI21X1 AOI21X1_219 ( .gnd(gnd), .vdd(vdd), .A(_2379_), .B(_2370_), .C(_2377_), .Y(_2383_) );
OAI21X1 OAI21X1_1295 ( .gnd(gnd), .vdd(vdd), .A(_2382_), .B(_2367_), .C(_2383_), .Y(_2384_) );
NOR2X1 NOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(_2368_), .B(_2382_), .Y(_2385_) );
AOI21X1 AOI21X1_220 ( .gnd(gnd), .vdd(vdd), .A(_2348_), .B(_2385_), .C(_2384_), .Y(_2386_) );
AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(_2385_), .B(_2345_), .Y(_2387_) );
OAI21X1 OAI21X1_1296 ( .gnd(gnd), .vdd(vdd), .A(_2315_), .B(_2318_), .C(_2387_), .Y(_2388_) );
NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_2386_), .B(_2388_), .Y(_2389_) );
NOR2X1 NOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(_794_), .B(_1650_), .Y(_2390_) );
NOR2X1 NOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(b_reg_16_), .B(_3667__112_), .Y(_2391_) );
NOR2X1 NOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(_2391_), .B(_2390_), .Y(_2392_) );
XNOR2X1 XNOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .B(_2392_), .Y(_2393_) );
OAI21X1 OAI21X1_1297 ( .gnd(gnd), .vdd(vdd), .A(_3667__112_), .B(_3432__bF_buf9), .C(_2005__bF_buf0), .Y(_2394_) );
OAI21X1 OAI21X1_1298 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf11), .B(_2393_), .C(_2394_), .Y(_1__16_) );
NOR2X1 NOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(_846_), .B(_1653_), .Y(_2395_) );
NOR2X1 NOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(b_reg_17_), .B(_3667__113_), .Y(_2396_) );
NOR2X1 NOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(_2396_), .B(_2395_), .Y(_2397_) );
INVX1 INVX1_925 ( .gnd(gnd), .vdd(vdd), .A(_2389_), .Y(_2398_) );
INVX1 INVX1_926 ( .gnd(gnd), .vdd(vdd), .A(_2390_), .Y(_2399_) );
OAI21X1 OAI21X1_1299 ( .gnd(gnd), .vdd(vdd), .A(_2391_), .B(_2398_), .C(_2399_), .Y(_2400_) );
NOR2X1 NOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(_2400_), .Y(_2401_) );
NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(_2400_), .Y(_2402_) );
NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf0), .B(_2402_), .Y(_2403_) );
OAI22X1 OAI22X1_85 ( .gnd(gnd), .vdd(vdd), .A(_1653_), .B(_2006__bF_buf6), .C(_2401_), .D(_2403_), .Y(_1__17_) );
NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_2392_), .B(_2397_), .Y(_2404_) );
AOI21X1 AOI21X1_221 ( .gnd(gnd), .vdd(vdd), .A(_2397_), .B(_2390_), .C(_2395_), .Y(_2405_) );
OAI21X1 OAI21X1_1300 ( .gnd(gnd), .vdd(vdd), .A(_2404_), .B(_2398_), .C(_2405_), .Y(_2406_) );
NOR2X1 NOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_1656_), .Y(_2407_) );
NOR2X1 NOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(b_reg_18_), .B(_3667__114_), .Y(_2408_) );
NOR2X1 NOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(_2408_), .B(_2407_), .Y(_2409_) );
NOR2X1 NOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(_2406_), .Y(_2410_) );
NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2409_), .B(_2406_), .Y(_2411_) );
NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(_2411_), .Y(_2412_) );
OAI21X1 OAI21X1_1301 ( .gnd(gnd), .vdd(vdd), .A(_3667__114_), .B(_3432__bF_buf8), .C(_2005__bF_buf10), .Y(_2413_) );
OAI21X1 OAI21X1_1302 ( .gnd(gnd), .vdd(vdd), .A(_2410_), .B(_2412_), .C(_2413_), .Y(_1__18_) );
OAI21X1 OAI21X1_1303 ( .gnd(gnd), .vdd(vdd), .A(_909_), .B(_1656_), .C(_2411_), .Y(_2414_) );
XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(b_reg_19_), .B(_3667__115_), .Y(_2415_) );
XNOR2X1 XNOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(_2414_), .B(_2415_), .Y(_2416_) );
OAI21X1 OAI21X1_1304 ( .gnd(gnd), .vdd(vdd), .A(_3667__115_), .B(_3432__bF_buf7), .C(_2005__bF_buf9), .Y(_2417_) );
OAI21X1 OAI21X1_1305 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf8), .B(_2416_), .C(_2417_), .Y(_1__19_) );
NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(_2415_), .B(_2409_), .Y(_2418_) );
NOR2X1 NOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .B(_2405_), .Y(_2419_) );
OAI21X1 OAI21X1_1306 ( .gnd(gnd), .vdd(vdd), .A(b_reg_19_), .B(_3667__115_), .C(_2407_), .Y(_2420_) );
OAI21X1 OAI21X1_1307 ( .gnd(gnd), .vdd(vdd), .A(_955_), .B(_1659_), .C(_2420_), .Y(_2421_) );
NOR2X1 NOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(_2421_), .B(_2419_), .Y(_2422_) );
NOR2X1 NOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(_2418_), .B(_2404_), .Y(_2423_) );
NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2423_), .B(_2389_), .Y(_2424_) );
AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(_2424_), .B(_2422_), .Y(_2425_) );
NOR2X1 NOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(_1023_), .B(_1662_), .Y(_2426_) );
NOR2X1 NOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(b_reg_20_), .B(_3667__116_), .Y(_2427_) );
NOR2X1 NOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(_2427_), .B(_2426_), .Y(_2428_) );
INVX1 INVX1_927 ( .gnd(gnd), .vdd(vdd), .A(_2428_), .Y(_2429_) );
NOR2X1 NOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(_2429_), .B(_2425_), .Y(_2430_) );
INVX1 INVX1_928 ( .gnd(gnd), .vdd(vdd), .A(_2425_), .Y(_2431_) );
OAI21X1 OAI21X1_1308 ( .gnd(gnd), .vdd(vdd), .A(_2428_), .B(_2431_), .C(digest_valid_new_bF_buf7), .Y(_2432_) );
OAI22X1 OAI22X1_86 ( .gnd(gnd), .vdd(vdd), .A(_1662_), .B(_2006__bF_buf5), .C(_2430_), .D(_2432_), .Y(_1__20_) );
NOR2X1 NOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1665_), .Y(_2433_) );
NOR2X1 NOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(b_reg_21_), .B(_3667__117_), .Y(_2434_) );
NOR2X1 NOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .B(_2430_), .Y(_2435_) );
OAI21X1 OAI21X1_1309 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_2434_), .C(_2435_), .Y(_2436_) );
NOR2X1 NOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(_2434_), .B(_2433_), .Y(_2437_) );
OAI21X1 OAI21X1_1310 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .B(_2430_), .C(_2437_), .Y(_2438_) );
NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2438_), .B(_2436_), .Y(_2439_) );
OAI22X1 OAI22X1_87 ( .gnd(gnd), .vdd(vdd), .A(_1665_), .B(_2006__bF_buf4), .C(_2005__bF_buf7), .D(_2439_), .Y(_1__21_) );
OAI21X1 OAI21X1_1311 ( .gnd(gnd), .vdd(vdd), .A(_1083_), .B(_1665_), .C(_2438_), .Y(_2440_) );
NOR2X1 NOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1668_), .Y(_2441_) );
NOR2X1 NOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(b_reg_22_), .B(_3667__118_), .Y(_2442_) );
NOR2X1 NOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(_2442_), .B(_2441_), .Y(_2443_) );
NOR2X1 NOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2440_), .Y(_2444_) );
NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2440_), .Y(_2445_) );
NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf6), .B(_2445_), .Y(_2446_) );
OAI21X1 OAI21X1_1312 ( .gnd(gnd), .vdd(vdd), .A(_3667__118_), .B(_3432__bF_buf6), .C(_2005__bF_buf6), .Y(_2447_) );
OAI21X1 OAI21X1_1313 ( .gnd(gnd), .vdd(vdd), .A(_2444_), .B(_2446_), .C(_2447_), .Y(_1__22_) );
OAI21X1 OAI21X1_1314 ( .gnd(gnd), .vdd(vdd), .A(_1141_), .B(_1668_), .C(_2445_), .Y(_2448_) );
NOR2X1 NOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(_1197_), .B(_1671_), .Y(_2449_) );
NOR2X1 NOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(b_reg_23_), .B(_3667__119_), .Y(_2450_) );
NOR2X1 NOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(_2450_), .B(_2449_), .Y(_2451_) );
XNOR2X1 XNOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(_2448_), .B(_2451_), .Y(_2452_) );
OAI21X1 OAI21X1_1315 ( .gnd(gnd), .vdd(vdd), .A(_3667__119_), .B(_3432__bF_buf5), .C(_2005__bF_buf5), .Y(_2453_) );
OAI21X1 OAI21X1_1316 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf4), .B(_2452_), .C(_2453_), .Y(_1__23_) );
NOR2X1 NOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(_1266_), .B(_1674_), .Y(_2454_) );
NOR2X1 NOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(b_reg_24_), .B(_3667__120_), .Y(_2455_) );
NOR2X1 NOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(_2455_), .B(_2454_), .Y(_2456_) );
INVX1 INVX1_929 ( .gnd(gnd), .vdd(vdd), .A(_2426_), .Y(_2457_) );
NOR2X1 NOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(_2434_), .B(_2457_), .Y(_2458_) );
NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(_2443_), .B(_2451_), .Y(_2459_) );
INVX1 INVX1_930 ( .gnd(gnd), .vdd(vdd), .A(_2459_), .Y(_2460_) );
OAI21X1 OAI21X1_1317 ( .gnd(gnd), .vdd(vdd), .A(_2433_), .B(_2458_), .C(_2460_), .Y(_2461_) );
AOI21X1 AOI21X1_222 ( .gnd(gnd), .vdd(vdd), .A(_2451_), .B(_2441_), .C(_2449_), .Y(_2462_) );
AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(_2461_), .B(_2462_), .Y(_2463_) );
AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(_2428_), .B(_2437_), .Y(_2464_) );
NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2460_), .Y(_2465_) );
OAI21X1 OAI21X1_1318 ( .gnd(gnd), .vdd(vdd), .A(_2465_), .B(_2422_), .C(_2463_), .Y(_2466_) );
NAND3X1 NAND3X1_300 ( .gnd(gnd), .vdd(vdd), .A(_2464_), .B(_2460_), .C(_2423_), .Y(_2467_) );
NOR2X1 NOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(_2467_), .B(_2398_), .Y(_2468_) );
NOR2X1 NOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(_2466_), .B(_2468_), .Y(_2469_) );
INVX1 INVX1_931 ( .gnd(gnd), .vdd(vdd), .A(_2469_), .Y(_2470_) );
NOR2X1 NOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(_2456_), .B(_2470_), .Y(_2471_) );
INVX1 INVX1_932 ( .gnd(gnd), .vdd(vdd), .A(_2456_), .Y(_2472_) );
OAI21X1 OAI21X1_1319 ( .gnd(gnd), .vdd(vdd), .A(_2472_), .B(_2469_), .C(digest_valid_new_bF_buf5), .Y(_2473_) );
OAI21X1 OAI21X1_1320 ( .gnd(gnd), .vdd(vdd), .A(_3667__120_), .B(_3432__bF_buf4), .C(_2005__bF_buf3), .Y(_2474_) );
OAI21X1 OAI21X1_1321 ( .gnd(gnd), .vdd(vdd), .A(_2473_), .B(_2471_), .C(_2474_), .Y(_1__24_) );
AOI21X1 AOI21X1_223 ( .gnd(gnd), .vdd(vdd), .A(_2470_), .B(_2456_), .C(_2454_), .Y(_2475_) );
NOR2X1 NOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(_1307_), .B(_1677_), .Y(_2476_) );
NOR2X1 NOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(b_reg_25_), .B(_3667__121_), .Y(_2477_) );
NOR2X1 NOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(_2477_), .B(_2476_), .Y(_2478_) );
INVX1 INVX1_933 ( .gnd(gnd), .vdd(vdd), .A(_2478_), .Y(_2479_) );
XNOR2X1 XNOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(_2475_), .B(_2479_), .Y(_2480_) );
OAI21X1 OAI21X1_1322 ( .gnd(gnd), .vdd(vdd), .A(_3667__121_), .B(_3432__bF_buf3), .C(_2005__bF_buf2), .Y(_2481_) );
OAI21X1 OAI21X1_1323 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf1), .B(_2480_), .C(_2481_), .Y(_1__25_) );
NOR2X1 NOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(_2472_), .B(_2479_), .Y(_2482_) );
INVX1 INVX1_934 ( .gnd(gnd), .vdd(vdd), .A(_2482_), .Y(_2483_) );
AOI21X1 AOI21X1_224 ( .gnd(gnd), .vdd(vdd), .A(_2478_), .B(_2454_), .C(_2476_), .Y(_2484_) );
OAI21X1 OAI21X1_1324 ( .gnd(gnd), .vdd(vdd), .A(_2483_), .B(_2469_), .C(_2484_), .Y(_2485_) );
INVX1 INVX1_935 ( .gnd(gnd), .vdd(vdd), .A(_2485_), .Y(_2486_) );
NOR2X1 NOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(_1680_), .Y(_2487_) );
NOR2X1 NOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(b_reg_26_), .B(_3667__122_), .Y(_2488_) );
OAI21X1 OAI21X1_1325 ( .gnd(gnd), .vdd(vdd), .A(_2487_), .B(_2488_), .C(_2486_), .Y(_2489_) );
NOR2X1 NOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(_2488_), .B(_2487_), .Y(_2490_) );
NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_2490_), .B(_2485_), .Y(_2491_) );
NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_2491_), .B(_2489_), .Y(_2492_) );
OAI21X1 OAI21X1_1326 ( .gnd(gnd), .vdd(vdd), .A(_3667__122_), .B(_3432__bF_buf2), .C(_2005__bF_buf0), .Y(_2493_) );
OAI21X1 OAI21X1_1327 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf11), .B(_2492_), .C(_2493_), .Y(_1__26_) );
OAI21X1 OAI21X1_1328 ( .gnd(gnd), .vdd(vdd), .A(_1347_), .B(_1680_), .C(_2491_), .Y(_2494_) );
AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(b_reg_27_), .B(_3667__123_), .Y(_2495_) );
NOR2X1 NOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(b_reg_27_), .B(_3667__123_), .Y(_2496_) );
NOR2X1 NOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(_2496_), .B(_2495_), .Y(_2497_) );
XNOR2X1 XNOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(_2494_), .B(_2497_), .Y(_2498_) );
OAI21X1 OAI21X1_1329 ( .gnd(gnd), .vdd(vdd), .A(_3667__123_), .B(_3432__bF_buf1), .C(_2005__bF_buf10), .Y(_2499_) );
OAI21X1 OAI21X1_1330 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf9), .B(_2498_), .C(_2499_), .Y(_1__27_) );
AOI21X1 AOI21X1_225 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .B(_2487_), .C(_2495_), .Y(_2500_) );
NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(_2497_), .B(_2490_), .Y(_2501_) );
OAI21X1 OAI21X1_1331 ( .gnd(gnd), .vdd(vdd), .A(_2501_), .B(_2486_), .C(_2500_), .Y(_2502_) );
XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(b_reg_28_), .B(_3667__124_), .Y(_2503_) );
NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_2502_), .Y(_2504_) );
INVX1 INVX1_936 ( .gnd(gnd), .vdd(vdd), .A(_2504_), .Y(_2505_) );
OAI21X1 OAI21X1_1332 ( .gnd(gnd), .vdd(vdd), .A(_2503_), .B(_2502_), .C(digest_valid_new_bF_buf4), .Y(_2506_) );
OAI22X1 OAI22X1_88 ( .gnd(gnd), .vdd(vdd), .A(_1685_), .B(_2006__bF_buf3), .C(_2506_), .D(_2505_), .Y(_1__28_) );
NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(b_reg_28_), .B(_3667__124_), .Y(_2507_) );
AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(_2504_), .B(_2507_), .Y(_2508_) );
NOR2X1 NOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(_1472_), .B(_1688_), .Y(_2509_) );
NOR2X1 NOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(b_reg_29_), .B(_3667__125_), .Y(_2510_) );
NOR2X1 NOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(_2510_), .B(_2509_), .Y(_2511_) );
AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(_2508_), .B(_2511_), .Y(_2512_) );
NOR2X1 NOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .B(_2508_), .Y(_2513_) );
OAI21X1 OAI21X1_1333 ( .gnd(gnd), .vdd(vdd), .A(_2513_), .B(_2512_), .C(digest_valid_new_bF_buf3), .Y(_2514_) );
OAI21X1 OAI21X1_1334 ( .gnd(gnd), .vdd(vdd), .A(_3667__125_), .B(_3432__bF_buf0), .C(_2005__bF_buf8), .Y(_2515_) );
NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_2515_), .B(_2514_), .Y(_1768_) );
XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(b_reg_30_), .B(_3667__126_), .Y(_2516_) );
INVX1 INVX1_937 ( .gnd(gnd), .vdd(vdd), .A(_2516_), .Y(_2517_) );
INVX1 INVX1_938 ( .gnd(gnd), .vdd(vdd), .A(_2509_), .Y(_2518_) );
OAI21X1 OAI21X1_1335 ( .gnd(gnd), .vdd(vdd), .A(_2507_), .B(_2510_), .C(_2518_), .Y(_2519_) );
AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(_2511_), .B(_2503_), .Y(_2520_) );
AOI21X1 AOI21X1_226 ( .gnd(gnd), .vdd(vdd), .A(_2502_), .B(_2520_), .C(_2519_), .Y(_2521_) );
AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(_2521_), .B(_2517_), .Y(_2522_) );
OAI21X1 OAI21X1_1336 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .B(_2521_), .C(digest_valid_new_bF_buf2), .Y(_2523_) );
OAI21X1 OAI21X1_1337 ( .gnd(gnd), .vdd(vdd), .A(_3667__126_), .B(_3432__bF_buf11), .C(_2005__bF_buf7), .Y(_2524_) );
OAI21X1 OAI21X1_1338 ( .gnd(gnd), .vdd(vdd), .A(_2522_), .B(_2523_), .C(_2524_), .Y(_1__30_) );
NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(b_reg_30_), .B(_3667__126_), .Y(_2525_) );
OAI21X1 OAI21X1_1339 ( .gnd(gnd), .vdd(vdd), .A(_2517_), .B(_2521_), .C(_2525_), .Y(_2526_) );
XNOR2X1 XNOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(b_reg_31_), .B(_3667__127_), .Y(_2527_) );
NOR2X1 NOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(_2527_), .B(_2526_), .Y(_2528_) );
AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(_2526_), .B(_2527_), .Y(_2529_) );
OAI21X1 OAI21X1_1340 ( .gnd(gnd), .vdd(vdd), .A(_2528_), .B(_2529_), .C(digest_valid_new_bF_buf1), .Y(_2530_) );
OAI21X1 OAI21X1_1341 ( .gnd(gnd), .vdd(vdd), .A(_3667__127_), .B(_3432__bF_buf10), .C(_2005__bF_buf6), .Y(_2531_) );
NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(_2531_), .B(_2530_), .Y(_1__31_) );
XNOR2X1 XNOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(c_reg_0_), .B(_3667__64_), .Y(_2532_) );
OAI22X1 OAI22X1_89 ( .gnd(gnd), .vdd(vdd), .A(_1695_), .B(_2006__bF_buf2), .C(_2005__bF_buf5), .D(_2532_), .Y(_2__0_) );
NOR2X1 NOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(_3413_), .B(_1695_), .Y(_2533_) );
XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(c_reg_1_), .B(_3667__65_), .Y(_2534_) );
XNOR2X1 XNOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(_2534_), .B(_2533_), .Y(_2535_) );
NOR2X1 NOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf0), .B(_1699_), .Y(_2536_) );
AOI21X1 AOI21X1_227 ( .gnd(gnd), .vdd(vdd), .A(_2535_), .B(digest_valid_new_bF_buf8), .C(_2536_), .Y(_2__1_) );
NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_2533_), .B(_2534_), .Y(_2537_) );
OAI21X1 OAI21X1_1342 ( .gnd(gnd), .vdd(vdd), .A(_3439_), .B(_1698_), .C(_2537_), .Y(_2538_) );
NOR2X1 NOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(_1701_), .B(_1702_), .Y(_2539_) );
NOR2X1 NOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(c_reg_2_), .B(_3667__66_), .Y(_2540_) );
NOR2X1 NOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(_2540_), .B(_2539_), .Y(_2541_) );
XNOR2X1 XNOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(_2538_), .B(_2541_), .Y(_2542_) );
NOR2X1 NOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf7), .B(_1703_), .Y(_2543_) );
AOI21X1 AOI21X1_228 ( .gnd(gnd), .vdd(vdd), .A(_2542_), .B(digest_valid_new_bF_buf6), .C(_2543_), .Y(_2__2_) );
AOI21X1 AOI21X1_229 ( .gnd(gnd), .vdd(vdd), .A(_2538_), .B(_2541_), .C(_2539_), .Y(_2544_) );
NOR2X1 NOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(_3574_), .B(_1705_), .Y(_2545_) );
NOR2X1 NOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(c_reg_3_), .B(_3667__67_), .Y(_2546_) );
NOR2X1 NOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(_2546_), .B(_2545_), .Y(_2547_) );
XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_2544_), .B(_2547_), .Y(_2548_) );
OAI21X1 OAI21X1_1343 ( .gnd(gnd), .vdd(vdd), .A(_3667__67_), .B(_3432__bF_buf9), .C(_2005__bF_buf4), .Y(_2549_) );
OAI21X1 OAI21X1_1344 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf3), .B(_2548_), .C(_2549_), .Y(_2__3_) );
XOR2X1 XOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(c_reg_4_), .B(_3667__68_), .Y(_2550_) );
INVX1 INVX1_939 ( .gnd(gnd), .vdd(vdd), .A(_2545_), .Y(_2551_) );
OAI21X1 OAI21X1_1345 ( .gnd(gnd), .vdd(vdd), .A(_2546_), .B(_2544_), .C(_2551_), .Y(_2552_) );
XNOR2X1 XNOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(_2552_), .B(_2550_), .Y(_2553_) );
NOR2X1 NOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf5), .B(_1709_), .Y(_2554_) );
AOI21X1 AOI21X1_230 ( .gnd(gnd), .vdd(vdd), .A(_2553_), .B(digest_valid_new_bF_buf4), .C(_2554_), .Y(_2__4_) );
NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_2550_), .B(_2552_), .Y(_2555_) );
OAI21X1 OAI21X1_1346 ( .gnd(gnd), .vdd(vdd), .A(_3641_), .B(_1708_), .C(_2555_), .Y(_2556_) );
XOR2X1 XOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(c_reg_5_), .B(_3667__69_), .Y(_2557_) );
NOR2X1 NOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(_2557_), .B(_2556_), .Y(_2558_) );
NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(_2557_), .B(_2556_), .Y(_2559_) );
NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf3), .B(_2559_), .Y(_2560_) );
OAI21X1 OAI21X1_1347 ( .gnd(gnd), .vdd(vdd), .A(_3667__69_), .B(_3432__bF_buf8), .C(_2005__bF_buf2), .Y(_2561_) );
OAI21X1 OAI21X1_1348 ( .gnd(gnd), .vdd(vdd), .A(_2558_), .B(_2560_), .C(_2561_), .Y(_2__5_) );
OAI21X1 OAI21X1_1349 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_1711_), .C(_2559_), .Y(_2562_) );
NOR2X1 NOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(_1714_), .B(_1715_), .Y(_2563_) );
NOR2X1 NOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(c_reg_6_), .B(_3667__70_), .Y(_2564_) );
NOR2X1 NOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(_2564_), .B(_2563_), .Y(_2565_) );
NOR2X1 NOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(_2565_), .B(_2562_), .Y(_2566_) );
NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_2565_), .B(_2562_), .Y(_2567_) );
NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf2), .B(_2567_), .Y(_2568_) );
OAI21X1 OAI21X1_1350 ( .gnd(gnd), .vdd(vdd), .A(_3667__70_), .B(_3432__bF_buf7), .C(_2005__bF_buf1), .Y(_2569_) );
OAI21X1 OAI21X1_1351 ( .gnd(gnd), .vdd(vdd), .A(_2566_), .B(_2568_), .C(_2569_), .Y(_2__6_) );
NOR2X1 NOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf1), .B(_1719_), .Y(_2570_) );
OAI21X1 OAI21X1_1352 ( .gnd(gnd), .vdd(vdd), .A(_1714_), .B(_1715_), .C(_2567_), .Y(_2571_) );
INVX1 INVX1_940 ( .gnd(gnd), .vdd(vdd), .A(_2571_), .Y(_2572_) );
NOR2X1 NOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(_189_), .B(_1718_), .Y(_2573_) );
NOR2X1 NOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(c_reg_7_), .B(_3667__71_), .Y(_2574_) );
NOR2X1 NOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .B(_2573_), .Y(_2575_) );
NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(_2575_), .B(_2572_), .Y(_2576_) );
NOR2X1 NOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(_2575_), .B(_2572_), .Y(_2577_) );
NOR2X1 NOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf0), .B(_2577_), .Y(_2578_) );
AOI21X1 AOI21X1_231 ( .gnd(gnd), .vdd(vdd), .A(_2578_), .B(_2576_), .C(_2570_), .Y(_2__7_) );
NOR2X1 NOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(_254_), .B(_1721_), .Y(_2579_) );
NOR2X1 NOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(c_reg_8_), .B(_3667__72_), .Y(_2580_) );
NOR2X1 NOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(_2580_), .B(_2579_), .Y(_2581_) );
INVX1 INVX1_941 ( .gnd(gnd), .vdd(vdd), .A(_2581_), .Y(_2582_) );
INVX1 INVX1_942 ( .gnd(gnd), .vdd(vdd), .A(_2574_), .Y(_2583_) );
OAI21X1 OAI21X1_1353 ( .gnd(gnd), .vdd(vdd), .A(_2573_), .B(_2571_), .C(_2583_), .Y(_2584_) );
NOR2X1 NOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(_2582_), .B(_2584_), .Y(_2585_) );
INVX1 INVX1_943 ( .gnd(gnd), .vdd(vdd), .A(_2584_), .Y(_2586_) );
OAI21X1 OAI21X1_1354 ( .gnd(gnd), .vdd(vdd), .A(_2581_), .B(_2586_), .C(digest_valid_new_bF_buf0), .Y(_2587_) );
OAI22X1 OAI22X1_90 ( .gnd(gnd), .vdd(vdd), .A(_1721_), .B(_2006__bF_buf1), .C(_2585_), .D(_2587_), .Y(_2__8_) );
NOR2X1 NOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_1724_), .Y(_2588_) );
NOR2X1 NOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(c_reg_9_), .B(_3667__73_), .Y(_2589_) );
NOR2X1 NOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .B(_2588_), .Y(_2590_) );
INVX1 INVX1_944 ( .gnd(gnd), .vdd(vdd), .A(_2579_), .Y(_2591_) );
OAI21X1 OAI21X1_1355 ( .gnd(gnd), .vdd(vdd), .A(_2580_), .B(_2584_), .C(_2591_), .Y(_2592_) );
NOR2X1 NOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(_2590_), .B(_2592_), .Y(_2593_) );
OAI21X1 OAI21X1_1356 ( .gnd(gnd), .vdd(vdd), .A(_2579_), .B(_2585_), .C(_2590_), .Y(_2594_) );
NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(_2594_), .Y(_2595_) );
OAI22X1 OAI22X1_91 ( .gnd(gnd), .vdd(vdd), .A(_1724_), .B(_2006__bF_buf0), .C(_2593_), .D(_2595_), .Y(_2__9_) );
OAI21X1 OAI21X1_1357 ( .gnd(gnd), .vdd(vdd), .A(_312_), .B(_1724_), .C(_2594_), .Y(_2596_) );
NOR2X1 NOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_1727_), .Y(_2597_) );
NOR2X1 NOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(c_reg_10_), .B(_3667__74_), .Y(_2598_) );
NOR2X1 NOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(_2598_), .B(_2597_), .Y(_2599_) );
NOR2X1 NOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(_2599_), .B(_2596_), .Y(_2600_) );
NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_2599_), .B(_2596_), .Y(_2601_) );
NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf7), .B(_2601_), .Y(_2602_) );
OAI21X1 OAI21X1_1358 ( .gnd(gnd), .vdd(vdd), .A(_3667__74_), .B(_3432__bF_buf6), .C(_2005__bF_buf11), .Y(_2603_) );
OAI21X1 OAI21X1_1359 ( .gnd(gnd), .vdd(vdd), .A(_2600_), .B(_2602_), .C(_2603_), .Y(_2__10_) );
OAI21X1 OAI21X1_1360 ( .gnd(gnd), .vdd(vdd), .A(_389_), .B(_1727_), .C(_2601_), .Y(_2604_) );
NOR2X1 NOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(_457_), .B(_1730_), .Y(_2605_) );
NOR2X1 NOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(c_reg_11_), .B(_3667__75_), .Y(_2606_) );
NOR2X1 NOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(_2606_), .B(_2605_), .Y(_2607_) );
XNOR2X1 XNOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(_2604_), .B(_2607_), .Y(_2608_) );
OAI21X1 OAI21X1_1361 ( .gnd(gnd), .vdd(vdd), .A(_3667__75_), .B(_3432__bF_buf5), .C(_2005__bF_buf10), .Y(_2609_) );
OAI21X1 OAI21X1_1362 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf9), .B(_2608_), .C(_2609_), .Y(_2__11_) );
AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(_2581_), .B(_2590_), .Y(_2610_) );
NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_2599_), .B(_2607_), .Y(_2611_) );
INVX1 INVX1_945 ( .gnd(gnd), .vdd(vdd), .A(_2611_), .Y(_2612_) );
NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(_2610_), .B(_2612_), .Y(_2613_) );
NOR2X1 NOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(_2589_), .B(_2591_), .Y(_2614_) );
OAI21X1 OAI21X1_1363 ( .gnd(gnd), .vdd(vdd), .A(_2588_), .B(_2614_), .C(_2612_), .Y(_2615_) );
AOI21X1 AOI21X1_232 ( .gnd(gnd), .vdd(vdd), .A(_2607_), .B(_2597_), .C(_2605_), .Y(_2616_) );
NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(_2616_), .B(_2615_), .Y(_2617_) );
INVX1 INVX1_946 ( .gnd(gnd), .vdd(vdd), .A(_2617_), .Y(_2618_) );
OAI21X1 OAI21X1_1364 ( .gnd(gnd), .vdd(vdd), .A(_2613_), .B(_2584_), .C(_2618_), .Y(_2619_) );
NOR2X1 NOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(_526_), .B(_1733_), .Y(_2620_) );
NOR2X1 NOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(c_reg_12_), .B(_3667__76_), .Y(_2621_) );
NOR2X1 NOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(_2621_), .B(_2620_), .Y(_2622_) );
NOR2X1 NOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(_2622_), .B(_2619_), .Y(_2623_) );
NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_2622_), .B(_2619_), .Y(_2624_) );
NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf6), .B(_2624_), .Y(_2625_) );
OAI21X1 OAI21X1_1365 ( .gnd(gnd), .vdd(vdd), .A(_3667__76_), .B(_3432__bF_buf4), .C(_2005__bF_buf8), .Y(_2626_) );
OAI21X1 OAI21X1_1366 ( .gnd(gnd), .vdd(vdd), .A(_2623_), .B(_2625_), .C(_2626_), .Y(_2__12_) );
INVX1 INVX1_947 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .Y(_2627_) );
NOR2X1 NOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(_588_), .B(_1736_), .Y(_2628_) );
NOR2X1 NOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(c_reg_13_), .B(_3667__77_), .Y(_2629_) );
NOR2X1 NOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(_2629_), .B(_2628_), .Y(_2630_) );
INVX1 INVX1_948 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .Y(_2631_) );
NAND3X1 NAND3X1_301 ( .gnd(gnd), .vdd(vdd), .A(_2627_), .B(_2631_), .C(_2624_), .Y(_2632_) );
NOR2X1 NOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(_2631_), .B(_2624_), .Y(_2633_) );
AOI21X1 AOI21X1_233 ( .gnd(gnd), .vdd(vdd), .A(_2620_), .B(_2630_), .C(_2633_), .Y(_2634_) );
NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_2632_), .B(_2634_), .Y(_2635_) );
OAI22X1 OAI22X1_92 ( .gnd(gnd), .vdd(vdd), .A(_1736_), .B(_2006__bF_buf8), .C(_2005__bF_buf7), .D(_2635_), .Y(_2__13_) );
AOI21X1 AOI21X1_234 ( .gnd(gnd), .vdd(vdd), .A(_2630_), .B(_2620_), .C(_2628_), .Y(_2636_) );
OAI21X1 OAI21X1_1367 ( .gnd(gnd), .vdd(vdd), .A(_2631_), .B(_2624_), .C(_2636_), .Y(_2637_) );
NOR2X1 NOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_1740_), .Y(_2638_) );
NOR2X1 NOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(c_reg_14_), .B(_3667__78_), .Y(_2639_) );
NOR2X1 NOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(_2639_), .B(_2638_), .Y(_2640_) );
NOR2X1 NOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(_2640_), .B(_2637_), .Y(_2641_) );
NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_2640_), .B(_2637_), .Y(_2642_) );
NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf5), .B(_2642_), .Y(_2643_) );
OAI21X1 OAI21X1_1368 ( .gnd(gnd), .vdd(vdd), .A(_3667__78_), .B(_3432__bF_buf3), .C(_2005__bF_buf6), .Y(_2644_) );
OAI21X1 OAI21X1_1369 ( .gnd(gnd), .vdd(vdd), .A(_2641_), .B(_2643_), .C(_2644_), .Y(_2__14_) );
OAI21X1 OAI21X1_1370 ( .gnd(gnd), .vdd(vdd), .A(_1739_), .B(_1740_), .C(_2642_), .Y(_2645_) );
NOR2X1 NOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(_744_), .B(_1743_), .Y(_2646_) );
NOR2X1 NOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(c_reg_15_), .B(_3667__79_), .Y(_2647_) );
NOR2X1 NOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(_2647_), .B(_2646_), .Y(_2648_) );
XNOR2X1 XNOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(_2645_), .B(_2648_), .Y(_2649_) );
OAI21X1 OAI21X1_1371 ( .gnd(gnd), .vdd(vdd), .A(_3667__79_), .B(_3432__bF_buf2), .C(_2005__bF_buf5), .Y(_2650_) );
OAI21X1 OAI21X1_1372 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf4), .B(_2649_), .C(_2650_), .Y(_2__15_) );
NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_2640_), .B(_2648_), .Y(_2651_) );
AOI21X1 AOI21X1_235 ( .gnd(gnd), .vdd(vdd), .A(_2648_), .B(_2638_), .C(_2646_), .Y(_2652_) );
OAI21X1 OAI21X1_1373 ( .gnd(gnd), .vdd(vdd), .A(_2651_), .B(_2636_), .C(_2652_), .Y(_2653_) );
NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_2622_), .B(_2630_), .Y(_2654_) );
NOR2X1 NOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(_2654_), .B(_2651_), .Y(_2655_) );
AOI21X1 AOI21X1_236 ( .gnd(gnd), .vdd(vdd), .A(_2617_), .B(_2655_), .C(_2653_), .Y(_2656_) );
NAND3X1 NAND3X1_302 ( .gnd(gnd), .vdd(vdd), .A(_2610_), .B(_2612_), .C(_2655_), .Y(_2657_) );
OAI21X1 OAI21X1_1374 ( .gnd(gnd), .vdd(vdd), .A(_2657_), .B(_2584_), .C(_2656_), .Y(_2658_) );
NOR2X1 NOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(_793_), .B(_1746_), .Y(_2659_) );
NOR2X1 NOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(c_reg_16_), .B(_3667__80_), .Y(_2660_) );
NOR2X1 NOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(_2660_), .B(_2659_), .Y(_2661_) );
AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2661_), .Y(_2662_) );
OAI21X1 OAI21X1_1375 ( .gnd(gnd), .vdd(vdd), .A(_2661_), .B(_2658_), .C(digest_valid_new_bF_buf4), .Y(_2663_) );
OAI22X1 OAI22X1_93 ( .gnd(gnd), .vdd(vdd), .A(_1746_), .B(_2006__bF_buf7), .C(_2662_), .D(_2663_), .Y(_2__16_) );
INVX1 INVX1_949 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .Y(_2664_) );
INVX1 INVX1_950 ( .gnd(gnd), .vdd(vdd), .A(_2659_), .Y(_2665_) );
OAI21X1 OAI21X1_1376 ( .gnd(gnd), .vdd(vdd), .A(_2660_), .B(_2664_), .C(_2665_), .Y(_2666_) );
NOR2X1 NOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_1749_), .Y(_2667_) );
NOR2X1 NOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(c_reg_17_), .B(_3667__81_), .Y(_2668_) );
NOR2X1 NOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(_2668_), .B(_2667_), .Y(_2669_) );
XNOR2X1 XNOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(_2666_), .B(_2669_), .Y(_2670_) );
OAI21X1 OAI21X1_1377 ( .gnd(gnd), .vdd(vdd), .A(_3667__81_), .B(_3432__bF_buf1), .C(_2005__bF_buf3), .Y(_2671_) );
OAI21X1 OAI21X1_1378 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf2), .B(_2670_), .C(_2671_), .Y(_2__17_) );
NOR2X1 NOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(_908_), .B(_1752_), .Y(_2672_) );
NOR2X1 NOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(c_reg_18_), .B(_3667__82_), .Y(_2673_) );
NOR2X1 NOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(_2673_), .B(_2672_), .Y(_2674_) );
INVX2 INVX2_83 ( .gnd(gnd), .vdd(vdd), .A(_2674_), .Y(_2675_) );
INVX1 INVX1_951 ( .gnd(gnd), .vdd(vdd), .A(_2668_), .Y(_2676_) );
OAI21X1 OAI21X1_1379 ( .gnd(gnd), .vdd(vdd), .A(_847_), .B(_1749_), .C(_2665_), .Y(_2677_) );
OAI21X1 OAI21X1_1380 ( .gnd(gnd), .vdd(vdd), .A(_2677_), .B(_2662_), .C(_2676_), .Y(_2678_) );
XNOR2X1 XNOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(_2678_), .B(_2675_), .Y(_2679_) );
OAI22X1 OAI22X1_94 ( .gnd(gnd), .vdd(vdd), .A(_1752_), .B(_2006__bF_buf6), .C(_2005__bF_buf1), .D(_2679_), .Y(_2__18_) );
INVX1 INVX1_952 ( .gnd(gnd), .vdd(vdd), .A(_2672_), .Y(_2680_) );
OAI21X1 OAI21X1_1381 ( .gnd(gnd), .vdd(vdd), .A(_2675_), .B(_2678_), .C(_2680_), .Y(_2681_) );
NOR2X1 NOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(_954_), .B(_1755_), .Y(_2682_) );
NOR2X1 NOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(c_reg_19_), .B(_3667__83_), .Y(_2683_) );
NOR2X1 NOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(_2683_), .B(_2682_), .Y(_2684_) );
INVX1 INVX1_953 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .Y(_2685_) );
NOR2X1 NOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(_2685_), .B(_2681_), .Y(_2686_) );
AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(_2681_), .B(_2685_), .Y(_2687_) );
OAI21X1 OAI21X1_1382 ( .gnd(gnd), .vdd(vdd), .A(_2686_), .B(_2687_), .C(digest_valid_new_bF_buf3), .Y(_2688_) );
OAI21X1 OAI21X1_1383 ( .gnd(gnd), .vdd(vdd), .A(_3667__83_), .B(_3432__bF_buf0), .C(_2005__bF_buf0), .Y(_2689_) );
NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(_2689_), .B(_2688_), .Y(_2__19_) );
OAI21X1 OAI21X1_1384 ( .gnd(gnd), .vdd(vdd), .A(c_reg_17_), .B(_3667__81_), .C(_2677_), .Y(_2690_) );
NOR2X1 NOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(_2675_), .B(_2685_), .Y(_2691_) );
INVX1 INVX1_954 ( .gnd(gnd), .vdd(vdd), .A(_2691_), .Y(_2692_) );
AOI21X1 AOI21X1_237 ( .gnd(gnd), .vdd(vdd), .A(_2684_), .B(_2672_), .C(_2682_), .Y(_2693_) );
OAI21X1 OAI21X1_1385 ( .gnd(gnd), .vdd(vdd), .A(_2690_), .B(_2692_), .C(_2693_), .Y(_2694_) );
NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_2661_), .B(_2669_), .Y(_2695_) );
NOR2X1 NOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(_2695_), .B(_2692_), .Y(_2696_) );
AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2696_), .Y(_2697_) );
NOR2X1 NOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .B(_2697_), .Y(_2698_) );
NOR2X1 NOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(_1022_), .B(_1758_), .Y(_2699_) );
NOR2X1 NOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(c_reg_20_), .B(_3667__84_), .Y(_2700_) );
OAI21X1 OAI21X1_1386 ( .gnd(gnd), .vdd(vdd), .A(_2699_), .B(_2700_), .C(_2698_), .Y(_2701_) );
NOR2X1 NOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(_2700_), .B(_2699_), .Y(_2702_) );
OAI21X1 OAI21X1_1387 ( .gnd(gnd), .vdd(vdd), .A(_2694_), .B(_2697_), .C(_2702_), .Y(_2703_) );
NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(_2703_), .B(_2701_), .Y(_2704_) );
OAI21X1 OAI21X1_1388 ( .gnd(gnd), .vdd(vdd), .A(_3667__84_), .B(_3432__bF_buf11), .C(_2005__bF_buf11), .Y(_2705_) );
OAI21X1 OAI21X1_1389 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf10), .B(_2704_), .C(_2705_), .Y(_2__20_) );
OAI21X1 OAI21X1_1390 ( .gnd(gnd), .vdd(vdd), .A(_1022_), .B(_1758_), .C(_2703_), .Y(_2706_) );
XOR2X1 XOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(c_reg_21_), .B(_3667__85_), .Y(_2707_) );
XNOR2X1 XNOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(_2706_), .B(_2707_), .Y(_2708_) );
OAI21X1 OAI21X1_1391 ( .gnd(gnd), .vdd(vdd), .A(_3667__85_), .B(_3432__bF_buf10), .C(_2005__bF_buf9), .Y(_2709_) );
OAI21X1 OAI21X1_1392 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf8), .B(_2708_), .C(_2709_), .Y(_2__21_) );
NOR2X1 NOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(_1140_), .B(_1764_), .Y(_2710_) );
NOR2X1 NOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(c_reg_22_), .B(_3667__86_), .Y(_2711_) );
NOR2X1 NOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(_2711_), .B(_2710_), .Y(_2712_) );
NOR2X1 NOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(_1082_), .B(_1761_), .Y(_2713_) );
AOI21X1 AOI21X1_238 ( .gnd(gnd), .vdd(vdd), .A(_2707_), .B(_2699_), .C(_2713_), .Y(_2714_) );
NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_2707_), .B(_2702_), .Y(_2715_) );
OAI21X1 OAI21X1_1393 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .B(_2698_), .C(_2714_), .Y(_2716_) );
AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(_2716_), .B(_2712_), .Y(_2717_) );
OAI21X1 OAI21X1_1394 ( .gnd(gnd), .vdd(vdd), .A(_2712_), .B(_2716_), .C(digest_valid_new_bF_buf2), .Y(_2718_) );
OAI22X1 OAI22X1_95 ( .gnd(gnd), .vdd(vdd), .A(_1764_), .B(_2006__bF_buf5), .C(_2717_), .D(_2718_), .Y(_2__22_) );
AOI21X1 AOI21X1_239 ( .gnd(gnd), .vdd(vdd), .A(_2716_), .B(_2712_), .C(_2710_), .Y(_2719_) );
NOR2X1 NOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(_1198_), .B(_1767_), .Y(_2720_) );
NOR2X1 NOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(c_reg_23_), .B(_3667__87_), .Y(_2721_) );
NOR2X1 NOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(_2721_), .B(_2720_), .Y(_2722_) );
XOR2X1 XOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_2719_), .B(_2722_), .Y(_2723_) );
OAI21X1 OAI21X1_1395 ( .gnd(gnd), .vdd(vdd), .A(_3667__87_), .B(_3432__bF_buf9), .C(_2005__bF_buf7), .Y(_2724_) );
OAI21X1 OAI21X1_1396 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf6), .B(_2723_), .C(_2724_), .Y(_2__23_) );
NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(_2712_), .B(_2722_), .Y(_2725_) );
NOR2X1 NOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(_2715_), .B(_2725_), .Y(_2726_) );
NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_2726_), .B(_2694_), .Y(_2727_) );
INVX1 INVX1_955 ( .gnd(gnd), .vdd(vdd), .A(_2727_), .Y(_2728_) );
AOI21X1 AOI21X1_240 ( .gnd(gnd), .vdd(vdd), .A(_2722_), .B(_2710_), .C(_2720_), .Y(_2729_) );
OAI21X1 OAI21X1_1397 ( .gnd(gnd), .vdd(vdd), .A(_2725_), .B(_2714_), .C(_2729_), .Y(_2730_) );
NOR2X1 NOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(_2730_), .B(_2728_), .Y(_2731_) );
INVX1 INVX1_956 ( .gnd(gnd), .vdd(vdd), .A(_2731_), .Y(_2732_) );
AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(_2696_), .B(_2726_), .Y(_2733_) );
AOI21X1 AOI21X1_241 ( .gnd(gnd), .vdd(vdd), .A(_2658_), .B(_2733_), .C(_2732_), .Y(_2734_) );
INVX1 INVX1_957 ( .gnd(gnd), .vdd(vdd), .A(_2734_), .Y(_2735_) );
NOR2X1 NOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(_1267_), .B(_1771_), .Y(_2736_) );
NOR2X1 NOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(c_reg_24_), .B(_3667__88_), .Y(_2737_) );
NOR2X1 NOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(_2737_), .B(_2736_), .Y(_2738_) );
AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(_2735_), .B(_2738_), .Y(_2739_) );
OAI21X1 OAI21X1_1398 ( .gnd(gnd), .vdd(vdd), .A(_2738_), .B(_2735_), .C(digest_valid_new_bF_buf1), .Y(_2740_) );
OAI22X1 OAI22X1_96 ( .gnd(gnd), .vdd(vdd), .A(_1771_), .B(_2006__bF_buf4), .C(_2739_), .D(_2740_), .Y(_2__24_) );
INVX1 INVX1_958 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .Y(_2741_) );
NOR2X1 NOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(_1308_), .B(_1774_), .Y(_2742_) );
NOR2X1 NOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(c_reg_25_), .B(_3667__89_), .Y(_2743_) );
OAI21X1 OAI21X1_1399 ( .gnd(gnd), .vdd(vdd), .A(_2742_), .B(_2743_), .C(_2741_), .Y(_2744_) );
NOR2X1 NOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(_2743_), .B(_2742_), .Y(_2745_) );
OAI21X1 OAI21X1_1400 ( .gnd(gnd), .vdd(vdd), .A(_2736_), .B(_2739_), .C(_2745_), .Y(_2746_) );
OAI21X1 OAI21X1_1401 ( .gnd(gnd), .vdd(vdd), .A(_2739_), .B(_2744_), .C(_2746_), .Y(_2747_) );
OAI22X1 OAI22X1_97 ( .gnd(gnd), .vdd(vdd), .A(_1774_), .B(_2006__bF_buf3), .C(_2005__bF_buf5), .D(_2747_), .Y(_2__25_) );
NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_2738_), .B(_2745_), .Y(_2748_) );
AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(_2745_), .B(_2736_), .Y(_2749_) );
NOR2X1 NOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(_2742_), .B(_2749_), .Y(_2750_) );
OAI21X1 OAI21X1_1402 ( .gnd(gnd), .vdd(vdd), .A(_2748_), .B(_2734_), .C(_2750_), .Y(_2751_) );
NOR2X1 NOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_1777_), .Y(_2752_) );
NOR2X1 NOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(c_reg_26_), .B(_3667__90_), .Y(_2753_) );
NOR2X1 NOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(_2753_), .B(_2752_), .Y(_2754_) );
NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_2751_), .Y(_2755_) );
INVX1 INVX1_959 ( .gnd(gnd), .vdd(vdd), .A(_2755_), .Y(_2756_) );
OAI21X1 OAI21X1_1403 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_2751_), .C(digest_valid_new_bF_buf0), .Y(_2757_) );
OAI22X1 OAI22X1_98 ( .gnd(gnd), .vdd(vdd), .A(_1777_), .B(_2006__bF_buf2), .C(_2757_), .D(_2756_), .Y(_2__26_) );
OAI21X1 OAI21X1_1404 ( .gnd(gnd), .vdd(vdd), .A(_1346_), .B(_1777_), .C(_2755_), .Y(_2758_) );
XOR2X1 XOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(c_reg_27_), .B(_3667__91_), .Y(_2759_) );
XNOR2X1 XNOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(_2758_), .B(_2759_), .Y(_2760_) );
OAI21X1 OAI21X1_1405 ( .gnd(gnd), .vdd(vdd), .A(_3667__91_), .B(_3432__bF_buf8), .C(_2005__bF_buf4), .Y(_2761_) );
OAI21X1 OAI21X1_1406 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf3), .B(_2760_), .C(_2761_), .Y(_2__27_) );
INVX1 INVX1_960 ( .gnd(gnd), .vdd(vdd), .A(_2750_), .Y(_2762_) );
OAI21X1 OAI21X1_1407 ( .gnd(gnd), .vdd(vdd), .A(c_reg_27_), .B(_3667__91_), .C(_2752_), .Y(_2763_) );
OAI21X1 OAI21X1_1408 ( .gnd(gnd), .vdd(vdd), .A(_1391_), .B(_1780_), .C(_2763_), .Y(_2764_) );
AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(_2754_), .B(_2759_), .Y(_2765_) );
AOI21X1 AOI21X1_242 ( .gnd(gnd), .vdd(vdd), .A(_2762_), .B(_2765_), .C(_2764_), .Y(_2766_) );
NAND3X1 NAND3X1_303 ( .gnd(gnd), .vdd(vdd), .A(_2738_), .B(_2745_), .C(_2765_), .Y(_2767_) );
OAI21X1 OAI21X1_1409 ( .gnd(gnd), .vdd(vdd), .A(_2767_), .B(_2734_), .C(_2766_), .Y(_2768_) );
NOR2X1 NOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1783_), .Y(_2769_) );
NOR2X1 NOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(c_reg_28_), .B(_3667__92_), .Y(_2770_) );
NOR2X1 NOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(_2770_), .B(_2769_), .Y(_2771_) );
NOR2X1 NOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(_2768_), .Y(_2772_) );
NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(_2768_), .Y(_2773_) );
NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(_2773_), .Y(_2774_) );
OAI21X1 OAI21X1_1410 ( .gnd(gnd), .vdd(vdd), .A(_3667__92_), .B(_3432__bF_buf7), .C(_2005__bF_buf2), .Y(_2775_) );
OAI21X1 OAI21X1_1411 ( .gnd(gnd), .vdd(vdd), .A(_2772_), .B(_2774_), .C(_2775_), .Y(_2__28_) );
OAI21X1 OAI21X1_1412 ( .gnd(gnd), .vdd(vdd), .A(_1434_), .B(_1783_), .C(_2773_), .Y(_2776_) );
NOR2X1 NOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(_1473_), .B(_1786_), .Y(_2777_) );
NOR2X1 NOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(c_reg_29_), .B(_3667__93_), .Y(_2778_) );
NOR2X1 NOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(_2778_), .B(_2777_), .Y(_2779_) );
AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(_2776_), .B(_2779_), .Y(_2780_) );
OAI21X1 OAI21X1_1413 ( .gnd(gnd), .vdd(vdd), .A(_2779_), .B(_2776_), .C(digest_valid_new_bF_buf7), .Y(_2781_) );
OAI22X1 OAI22X1_99 ( .gnd(gnd), .vdd(vdd), .A(_1786_), .B(_2006__bF_buf1), .C(_2780_), .D(_2781_), .Y(_2__29_) );
NOR2X1 NOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1789_), .Y(_2782_) );
INVX1 INVX1_961 ( .gnd(gnd), .vdd(vdd), .A(_2782_), .Y(_2783_) );
NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(_1524_), .B(_1789_), .Y(_2784_) );
AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(_2783_), .B(_2784_), .Y(_2785_) );
INVX1 INVX1_962 ( .gnd(gnd), .vdd(vdd), .A(_2785_), .Y(_2786_) );
INVX1 INVX1_963 ( .gnd(gnd), .vdd(vdd), .A(_2778_), .Y(_2787_) );
AOI21X1 AOI21X1_243 ( .gnd(gnd), .vdd(vdd), .A(_2769_), .B(_2787_), .C(_2777_), .Y(_2788_) );
INVX1 INVX1_964 ( .gnd(gnd), .vdd(vdd), .A(_2788_), .Y(_2789_) );
AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(_2771_), .B(_2779_), .Y(_2790_) );
AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(_2768_), .B(_2790_), .Y(_2791_) );
NOR2X1 NOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(_2789_), .B(_2791_), .Y(_2792_) );
AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(_2792_), .B(_2786_), .Y(_2793_) );
OAI21X1 OAI21X1_1414 ( .gnd(gnd), .vdd(vdd), .A(_2786_), .B(_2792_), .C(digest_valid_new_bF_buf6), .Y(_2794_) );
OAI22X1 OAI22X1_100 ( .gnd(gnd), .vdd(vdd), .A(_1789_), .B(_2006__bF_buf0), .C(_2793_), .D(_2794_), .Y(_2__30_) );
OAI21X1 OAI21X1_1415 ( .gnd(gnd), .vdd(vdd), .A(_2789_), .B(_2791_), .C(_2785_), .Y(_2795_) );
XNOR2X1 XNOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(c_reg_31_), .B(_3667__95_), .Y(_2796_) );
NAND3X1 NAND3X1_304 ( .gnd(gnd), .vdd(vdd), .A(_2783_), .B(_2796_), .C(_2795_), .Y(_2797_) );
NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_2790_), .B(_2768_), .Y(_2798_) );
AOI21X1 AOI21X1_244 ( .gnd(gnd), .vdd(vdd), .A(_2798_), .B(_2788_), .C(_2786_), .Y(_2799_) );
INVX1 INVX1_965 ( .gnd(gnd), .vdd(vdd), .A(_2796_), .Y(_2800_) );
OAI21X1 OAI21X1_1416 ( .gnd(gnd), .vdd(vdd), .A(_2782_), .B(_2799_), .C(_2800_), .Y(_2801_) );
NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_2801_), .B(_2797_), .Y(_2802_) );
OAI21X1 OAI21X1_1417 ( .gnd(gnd), .vdd(vdd), .A(_3667__95_), .B(_3432__bF_buf6), .C(_2005__bF_buf1), .Y(_2803_) );
OAI21X1 OAI21X1_1418 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf0), .B(_2802_), .C(_2803_), .Y(_2__31_) );
XNOR2X1 XNOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(d_reg_0_), .B(_3667__32_), .Y(_2804_) );
OAI22X1 OAI22X1_101 ( .gnd(gnd), .vdd(vdd), .A(_1794_), .B(_2006__bF_buf8), .C(_2005__bF_buf11), .D(_2804_), .Y(_3__0_) );
NOR2X1 NOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(_3393_), .B(_1794_), .Y(_2805_) );
XOR2X1 XOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(d_reg_1_), .B(_3667__33_), .Y(_2806_) );
XNOR2X1 XNOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(_2806_), .B(_2805_), .Y(_2807_) );
NOR2X1 NOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf5), .B(_1798_), .Y(_2808_) );
AOI21X1 AOI21X1_245 ( .gnd(gnd), .vdd(vdd), .A(_2807_), .B(digest_valid_new_bF_buf4), .C(_2808_), .Y(_3__1_) );
NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_2805_), .B(_2806_), .Y(_2809_) );
OAI21X1 OAI21X1_1419 ( .gnd(gnd), .vdd(vdd), .A(_3443_), .B(_1797_), .C(_2809_), .Y(_2810_) );
NOR2X1 NOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(_3508_), .B(_1800_), .Y(_2811_) );
NOR2X1 NOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(d_reg_2_), .B(_3667__34_), .Y(_2812_) );
NOR2X1 NOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(_2812_), .B(_2811_), .Y(_2813_) );
XNOR2X1 XNOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(_2810_), .B(_2813_), .Y(_2814_) );
NOR2X1 NOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf3), .B(_1801_), .Y(_2815_) );
AOI21X1 AOI21X1_246 ( .gnd(gnd), .vdd(vdd), .A(_2814_), .B(digest_valid_new_bF_buf2), .C(_2815_), .Y(_3__2_) );
AOI21X1 AOI21X1_247 ( .gnd(gnd), .vdd(vdd), .A(_2810_), .B(_2813_), .C(_2811_), .Y(_2816_) );
NOR2X1 NOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(_3573_), .B(_1803_), .Y(_2817_) );
NOR2X1 NOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(d_reg_3_), .B(_3667__35_), .Y(_2818_) );
NOR2X1 NOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(_2818_), .B(_2817_), .Y(_2819_) );
XOR2X1 XOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(_2816_), .B(_2819_), .Y(_2820_) );
OAI22X1 OAI22X1_102 ( .gnd(gnd), .vdd(vdd), .A(_1803_), .B(_2006__bF_buf7), .C(_2005__bF_buf10), .D(_2820_), .Y(_3__3_) );
XOR2X1 XOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(d_reg_4_), .B(_3667__36_), .Y(_2821_) );
INVX1 INVX1_966 ( .gnd(gnd), .vdd(vdd), .A(_2817_), .Y(_2822_) );
OAI21X1 OAI21X1_1420 ( .gnd(gnd), .vdd(vdd), .A(_2818_), .B(_2816_), .C(_2822_), .Y(_2823_) );
XNOR2X1 XNOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(_2823_), .B(_2821_), .Y(_2824_) );
NOR2X1 NOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf1), .B(_1807_), .Y(_2825_) );
AOI21X1 AOI21X1_248 ( .gnd(gnd), .vdd(vdd), .A(_2824_), .B(digest_valid_new_bF_buf0), .C(_2825_), .Y(_3__4_) );
NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_2821_), .B(_2823_), .Y(_2826_) );
OAI21X1 OAI21X1_1421 ( .gnd(gnd), .vdd(vdd), .A(_3639_), .B(_1806_), .C(_2826_), .Y(_2827_) );
XOR2X1 XOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(d_reg_5_), .B(_3667__37_), .Y(_2828_) );
NOR2X1 NOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(_2828_), .B(_2827_), .Y(_2829_) );
NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_2828_), .B(_2827_), .Y(_2830_) );
NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(_2830_), .Y(_2831_) );
OAI21X1 OAI21X1_1422 ( .gnd(gnd), .vdd(vdd), .A(_3667__37_), .B(_3432__bF_buf5), .C(_2005__bF_buf9), .Y(_2832_) );
OAI21X1 OAI21X1_1423 ( .gnd(gnd), .vdd(vdd), .A(_2829_), .B(_2831_), .C(_2832_), .Y(_3__5_) );
OAI21X1 OAI21X1_1424 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_1809_), .C(_2830_), .Y(_2833_) );
XOR2X1 XOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(d_reg_6_), .B(_3667__38_), .Y(_2834_) );
NOR2X1 NOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2833_), .Y(_2835_) );
NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_2834_), .B(_2833_), .Y(_2836_) );
NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf7), .B(_2836_), .Y(_2837_) );
OAI21X1 OAI21X1_1425 ( .gnd(gnd), .vdd(vdd), .A(_3667__38_), .B(_3432__bF_buf4), .C(_2005__bF_buf8), .Y(_2838_) );
OAI21X1 OAI21X1_1426 ( .gnd(gnd), .vdd(vdd), .A(_2835_), .B(_2837_), .C(_2838_), .Y(_3__6_) );
NOR2X1 NOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_1815_), .Y(_2839_) );
NOR2X1 NOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(d_reg_7_), .B(_3667__39_), .Y(_2840_) );
NOR2X1 NOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(_2840_), .B(_2839_), .Y(_2841_) );
OAI21X1 OAI21X1_1427 ( .gnd(gnd), .vdd(vdd), .A(_131_), .B(_1812_), .C(_2836_), .Y(_2842_) );
XNOR2X1 XNOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(_2842_), .B(_2841_), .Y(_2843_) );
OAI22X1 OAI22X1_103 ( .gnd(gnd), .vdd(vdd), .A(_1815_), .B(_2006__bF_buf6), .C(_2005__bF_buf7), .D(_2843_), .Y(_3__7_) );
AOI21X1 AOI21X1_249 ( .gnd(gnd), .vdd(vdd), .A(_2842_), .B(_2841_), .C(_2839_), .Y(_2844_) );
NOR2X1 NOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_1818_), .Y(_2845_) );
NOR2X1 NOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(d_reg_8_), .B(_3667__40_), .Y(_2846_) );
NOR2X1 NOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(_2846_), .B(_2845_), .Y(_2847_) );
INVX1 INVX1_967 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .Y(_2848_) );
NOR2X1 NOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(_2848_), .B(_2844_), .Y(_2849_) );
INVX1 INVX1_968 ( .gnd(gnd), .vdd(vdd), .A(_2844_), .Y(_2850_) );
OAI21X1 OAI21X1_1428 ( .gnd(gnd), .vdd(vdd), .A(_2847_), .B(_2850_), .C(digest_valid_new_bF_buf6), .Y(_2851_) );
OAI22X1 OAI22X1_104 ( .gnd(gnd), .vdd(vdd), .A(_1818_), .B(_2006__bF_buf5), .C(_2849_), .D(_2851_), .Y(_3__8_) );
NOR2X1 NOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(_310_), .B(_1821_), .Y(_2852_) );
NOR2X1 NOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(d_reg_9_), .B(_3667__41_), .Y(_2853_) );
NOR2X1 NOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(_2853_), .B(_2852_), .Y(_2854_) );
INVX1 INVX1_969 ( .gnd(gnd), .vdd(vdd), .A(_2854_), .Y(_2855_) );
NOR2X1 NOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(_2845_), .B(_2849_), .Y(_2856_) );
AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(_2856_), .B(_2855_), .Y(_2857_) );
OAI21X1 OAI21X1_1429 ( .gnd(gnd), .vdd(vdd), .A(_2855_), .B(_2856_), .C(digest_valid_new_bF_buf5), .Y(_2858_) );
OAI22X1 OAI22X1_105 ( .gnd(gnd), .vdd(vdd), .A(_1821_), .B(_2006__bF_buf4), .C(_2857_), .D(_2858_), .Y(_3__9_) );
NOR2X1 NOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(_2848_), .B(_2855_), .Y(_2859_) );
INVX1 INVX1_970 ( .gnd(gnd), .vdd(vdd), .A(_2859_), .Y(_2860_) );
AOI21X1 AOI21X1_250 ( .gnd(gnd), .vdd(vdd), .A(_2854_), .B(_2845_), .C(_2852_), .Y(_2861_) );
OAI21X1 OAI21X1_1430 ( .gnd(gnd), .vdd(vdd), .A(_2860_), .B(_2844_), .C(_2861_), .Y(_2862_) );
NOR2X1 NOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_1824_), .Y(_2863_) );
NOR2X1 NOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(d_reg_10_), .B(_3667__42_), .Y(_2864_) );
NOR2X1 NOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(_2864_), .B(_2863_), .Y(_2865_) );
NOR2X1 NOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(_2865_), .B(_2862_), .Y(_2866_) );
NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(_2865_), .B(_2862_), .Y(_2867_) );
NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf4), .B(_2867_), .Y(_2868_) );
OAI21X1 OAI21X1_1431 ( .gnd(gnd), .vdd(vdd), .A(_3667__42_), .B(_3432__bF_buf3), .C(_2005__bF_buf6), .Y(_2869_) );
OAI21X1 OAI21X1_1432 ( .gnd(gnd), .vdd(vdd), .A(_2866_), .B(_2868_), .C(_2869_), .Y(_3__10_) );
OAI21X1 OAI21X1_1433 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_1824_), .C(_2867_), .Y(_2870_) );
NOR2X1 NOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(_451_), .B(_1827_), .Y(_2871_) );
NOR2X1 NOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(d_reg_11_), .B(_3667__43_), .Y(_2872_) );
NOR2X1 NOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(_2872_), .B(_2871_), .Y(_2873_) );
XNOR2X1 XNOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(_2870_), .B(_2873_), .Y(_2874_) );
OAI22X1 OAI22X1_106 ( .gnd(gnd), .vdd(vdd), .A(_1827_), .B(_2006__bF_buf3), .C(_2005__bF_buf5), .D(_2874_), .Y(_3__11_) );
NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_2865_), .B(_2873_), .Y(_2875_) );
NOR2X1 NOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(_2875_), .B(_2860_), .Y(_2876_) );
INVX1 INVX1_971 ( .gnd(gnd), .vdd(vdd), .A(_2876_), .Y(_2877_) );
AOI21X1 AOI21X1_251 ( .gnd(gnd), .vdd(vdd), .A(_2873_), .B(_2863_), .C(_2871_), .Y(_2878_) );
OAI21X1 OAI21X1_1434 ( .gnd(gnd), .vdd(vdd), .A(_2875_), .B(_2861_), .C(_2878_), .Y(_2879_) );
INVX1 INVX1_972 ( .gnd(gnd), .vdd(vdd), .A(_2879_), .Y(_2880_) );
OAI21X1 OAI21X1_1435 ( .gnd(gnd), .vdd(vdd), .A(_2877_), .B(_2844_), .C(_2880_), .Y(_2881_) );
NOR2X1 NOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(_519_), .B(_1830_), .Y(_2882_) );
NOR2X1 NOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(d_reg_12_), .B(_3667__44_), .Y(_2883_) );
NOR2X1 NOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(_2883_), .B(_2882_), .Y(_2884_) );
AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_2884_), .Y(_2885_) );
NOR2X1 NOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf4), .B(_2885_), .Y(_2886_) );
OAI21X1 OAI21X1_1436 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_2884_), .C(_2886_), .Y(_2887_) );
OAI21X1 OAI21X1_1437 ( .gnd(gnd), .vdd(vdd), .A(_3667__44_), .B(_3432__bF_buf2), .C(_2005__bF_buf3), .Y(_2888_) );
NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_2888_), .B(_2887_), .Y(_3__12_) );
NOR2X1 NOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_1833_), .Y(_2889_) );
NOR2X1 NOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(d_reg_13_), .B(_3667__45_), .Y(_2890_) );
NOR2X1 NOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(_2882_), .B(_2885_), .Y(_2891_) );
OAI21X1 OAI21X1_1438 ( .gnd(gnd), .vdd(vdd), .A(_2889_), .B(_2890_), .C(_2891_), .Y(_2892_) );
NOR2X1 NOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(_2890_), .B(_2889_), .Y(_2893_) );
OAI21X1 OAI21X1_1439 ( .gnd(gnd), .vdd(vdd), .A(_2882_), .B(_2885_), .C(_2893_), .Y(_2894_) );
NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(_2894_), .B(_2892_), .Y(_2895_) );
OAI22X1 OAI22X1_107 ( .gnd(gnd), .vdd(vdd), .A(_1833_), .B(_2006__bF_buf2), .C(_2005__bF_buf2), .D(_2895_), .Y(_3__13_) );
AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(_2884_), .B(_2893_), .Y(_2896_) );
OAI21X1 OAI21X1_1440 ( .gnd(gnd), .vdd(vdd), .A(d_reg_13_), .B(_3667__45_), .C(_2882_), .Y(_2897_) );
OAI21X1 OAI21X1_1441 ( .gnd(gnd), .vdd(vdd), .A(_582_), .B(_1833_), .C(_2897_), .Y(_2898_) );
AOI21X1 AOI21X1_252 ( .gnd(gnd), .vdd(vdd), .A(_2881_), .B(_2896_), .C(_2898_), .Y(_2899_) );
NOR2X1 NOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(_653_), .B(_1836_), .Y(_2900_) );
NOR2X1 NOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(d_reg_14_), .B(_3667__46_), .Y(_2901_) );
NOR2X1 NOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(_2901_), .B(_2900_), .Y(_2902_) );
INVX2 INVX2_84 ( .gnd(gnd), .vdd(vdd), .A(_2902_), .Y(_2903_) );
AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(_2899_), .B(_2903_), .Y(_2904_) );
OAI21X1 OAI21X1_1442 ( .gnd(gnd), .vdd(vdd), .A(_2903_), .B(_2899_), .C(digest_valid_new_bF_buf3), .Y(_2905_) );
OAI21X1 OAI21X1_1443 ( .gnd(gnd), .vdd(vdd), .A(_3667__46_), .B(_3432__bF_buf1), .C(_2005__bF_buf1), .Y(_2906_) );
OAI21X1 OAI21X1_1444 ( .gnd(gnd), .vdd(vdd), .A(_2904_), .B(_2905_), .C(_2906_), .Y(_3__14_) );
INVX1 INVX1_973 ( .gnd(gnd), .vdd(vdd), .A(_2900_), .Y(_2907_) );
OAI21X1 OAI21X1_1445 ( .gnd(gnd), .vdd(vdd), .A(_2903_), .B(_2899_), .C(_2907_), .Y(_2908_) );
NOR2X1 NOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(_718_), .B(_1839_), .Y(_2909_) );
NOR2X1 NOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(d_reg_15_), .B(_3667__47_), .Y(_2910_) );
NOR2X1 NOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(_2910_), .B(_2909_), .Y(_2911_) );
INVX1 INVX1_974 ( .gnd(gnd), .vdd(vdd), .A(_2911_), .Y(_2912_) );
NOR2X1 NOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(_2912_), .B(_2908_), .Y(_2913_) );
AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(_2908_), .B(_2912_), .Y(_2914_) );
OAI21X1 OAI21X1_1446 ( .gnd(gnd), .vdd(vdd), .A(_2913_), .B(_2914_), .C(digest_valid_new_bF_buf2), .Y(_2915_) );
OAI21X1 OAI21X1_1447 ( .gnd(gnd), .vdd(vdd), .A(_1839_), .B(_2006__bF_buf1), .C(_2915_), .Y(_3__15_) );
NOR2X1 NOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(_2903_), .B(_2912_), .Y(_2916_) );
NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_2898_), .B(_2916_), .Y(_2917_) );
AOI21X1 AOI21X1_253 ( .gnd(gnd), .vdd(vdd), .A(_2911_), .B(_2900_), .C(_2909_), .Y(_2918_) );
NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_2918_), .B(_2917_), .Y(_2919_) );
AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(_2916_), .B(_2896_), .Y(_2920_) );
AOI21X1 AOI21X1_254 ( .gnd(gnd), .vdd(vdd), .A(_2879_), .B(_2920_), .C(_2919_), .Y(_2921_) );
NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(_2920_), .B(_2876_), .Y(_2922_) );
OAI21X1 OAI21X1_1448 ( .gnd(gnd), .vdd(vdd), .A(_2922_), .B(_2844_), .C(_2921_), .Y(_2923_) );
NOR2X1 NOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(_788_), .B(_1842_), .Y(_2924_) );
NOR2X1 NOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(d_reg_16_), .B(_3667__48_), .Y(_2925_) );
NOR2X1 NOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(_2925_), .B(_2924_), .Y(_2926_) );
AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(_2923_), .B(_2926_), .Y(_2927_) );
OAI21X1 OAI21X1_1449 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(_2923_), .C(digest_valid_new_bF_buf1), .Y(_2928_) );
OAI22X1 OAI22X1_108 ( .gnd(gnd), .vdd(vdd), .A(_1842_), .B(_2006__bF_buf0), .C(_2927_), .D(_2928_), .Y(_3__16_) );
NOR2X1 NOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_2927_), .Y(_2929_) );
NOR2X1 NOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(_853_), .B(_1845_), .Y(_2930_) );
NOR2X1 NOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(d_reg_17_), .B(_3667__49_), .Y(_2931_) );
NOR2X1 NOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(_2931_), .B(_2930_), .Y(_2932_) );
XOR2X1 XOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_2929_), .B(_2932_), .Y(_2933_) );
OAI21X1 OAI21X1_1450 ( .gnd(gnd), .vdd(vdd), .A(_3667__49_), .B(_3432__bF_buf0), .C(_2005__bF_buf0), .Y(_2934_) );
OAI21X1 OAI21X1_1451 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf11), .B(_2933_), .C(_2934_), .Y(_3__17_) );
NOR2X1 NOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(_903_), .B(_1848_), .Y(_2935_) );
NOR2X1 NOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(d_reg_18_), .B(_3667__50_), .Y(_2936_) );
NOR2X1 NOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(_2936_), .B(_2935_), .Y(_2937_) );
INVX1 INVX1_975 ( .gnd(gnd), .vdd(vdd), .A(_2937_), .Y(_2938_) );
INVX1 INVX1_976 ( .gnd(gnd), .vdd(vdd), .A(_2931_), .Y(_2939_) );
OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(_2924_), .B(_2930_), .Y(_2940_) );
OAI21X1 OAI21X1_1452 ( .gnd(gnd), .vdd(vdd), .A(_2940_), .B(_2927_), .C(_2939_), .Y(_2941_) );
NOR2X1 NOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(_2938_), .B(_2941_), .Y(_2942_) );
OAI21X1 OAI21X1_1453 ( .gnd(gnd), .vdd(vdd), .A(_2935_), .B(_2936_), .C(_2941_), .Y(_2943_) );
NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf0), .B(_2943_), .Y(_2944_) );
OAI22X1 OAI22X1_109 ( .gnd(gnd), .vdd(vdd), .A(_1848_), .B(_2006__bF_buf8), .C(_2942_), .D(_2944_), .Y(_3__18_) );
NOR2X1 NOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(_949_), .B(_1851_), .Y(_2945_) );
NOR2X1 NOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(d_reg_19_), .B(_3667__51_), .Y(_2946_) );
NOR2X1 NOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(_2946_), .B(_2945_), .Y(_2947_) );
OAI21X1 OAI21X1_1454 ( .gnd(gnd), .vdd(vdd), .A(_2935_), .B(_2942_), .C(_2947_), .Y(_2948_) );
NOR2X1 NOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(_2935_), .B(_2942_), .Y(_2949_) );
OAI21X1 OAI21X1_1455 ( .gnd(gnd), .vdd(vdd), .A(_2945_), .B(_2946_), .C(_2949_), .Y(_2950_) );
NAND3X1 NAND3X1_305 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(_2948_), .C(_2950_), .Y(_2951_) );
OAI21X1 OAI21X1_1456 ( .gnd(gnd), .vdd(vdd), .A(_1851_), .B(_2006__bF_buf7), .C(_2951_), .Y(_3__19_) );
OAI21X1 OAI21X1_1457 ( .gnd(gnd), .vdd(vdd), .A(d_reg_17_), .B(_3667__49_), .C(_2940_), .Y(_2952_) );
NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(_2937_), .B(_2947_), .Y(_2953_) );
AOI21X1 AOI21X1_255 ( .gnd(gnd), .vdd(vdd), .A(_2947_), .B(_2935_), .C(_2945_), .Y(_2954_) );
OAI21X1 OAI21X1_1458 ( .gnd(gnd), .vdd(vdd), .A(_2953_), .B(_2952_), .C(_2954_), .Y(_2955_) );
NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(_2926_), .B(_2932_), .Y(_2956_) );
NOR2X1 NOR2X1_563 ( .gnd(gnd), .vdd(vdd), .A(_2956_), .B(_2953_), .Y(_2957_) );
AOI21X1 AOI21X1_256 ( .gnd(gnd), .vdd(vdd), .A(_2923_), .B(_2957_), .C(_2955_), .Y(_2958_) );
NOR2X1 NOR2X1_564 ( .gnd(gnd), .vdd(vdd), .A(_1024_), .B(_1854_), .Y(_2959_) );
NOR2X1 NOR2X1_565 ( .gnd(gnd), .vdd(vdd), .A(d_reg_20_), .B(_3667__52_), .Y(_2960_) );
NOR2X1 NOR2X1_566 ( .gnd(gnd), .vdd(vdd), .A(_2960_), .B(_2959_), .Y(_2961_) );
INVX1 INVX1_977 ( .gnd(gnd), .vdd(vdd), .A(_2961_), .Y(_2962_) );
AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .B(_2962_), .Y(_2963_) );
OAI21X1 OAI21X1_1459 ( .gnd(gnd), .vdd(vdd), .A(_2962_), .B(_2958_), .C(digest_valid_new_bF_buf7), .Y(_2964_) );
OAI21X1 OAI21X1_1460 ( .gnd(gnd), .vdd(vdd), .A(_3667__52_), .B(_3432__bF_buf11), .C(_2005__bF_buf10), .Y(_2965_) );
OAI21X1 OAI21X1_1461 ( .gnd(gnd), .vdd(vdd), .A(_2963_), .B(_2964_), .C(_2965_), .Y(_3__20_) );
INVX1 INVX1_978 ( .gnd(gnd), .vdd(vdd), .A(_2958_), .Y(_2966_) );
AOI21X1 AOI21X1_257 ( .gnd(gnd), .vdd(vdd), .A(_2966_), .B(_2961_), .C(_2959_), .Y(_2967_) );
XOR2X1 XOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(d_reg_21_), .B(_3667__53_), .Y(_2968_) );
AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(_2967_), .B(_2968_), .Y(_2969_) );
NOR2X1 NOR2X1_567 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(_2967_), .Y(_2970_) );
OAI21X1 OAI21X1_1462 ( .gnd(gnd), .vdd(vdd), .A(_2970_), .B(_2969_), .C(digest_valid_new_bF_buf6), .Y(_2971_) );
OAI21X1 OAI21X1_1463 ( .gnd(gnd), .vdd(vdd), .A(_3667__53_), .B(_3432__bF_buf10), .C(_2005__bF_buf9), .Y(_2972_) );
NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_2972_), .B(_2971_), .Y(_3__21_) );
NOR2X1 NOR2X1_568 ( .gnd(gnd), .vdd(vdd), .A(_1142_), .B(_1860_), .Y(_2973_) );
NOR2X1 NOR2X1_569 ( .gnd(gnd), .vdd(vdd), .A(d_reg_22_), .B(_3667__54_), .Y(_2974_) );
NOR2X1 NOR2X1_570 ( .gnd(gnd), .vdd(vdd), .A(_2974_), .B(_2973_), .Y(_2975_) );
NOR2X1 NOR2X1_571 ( .gnd(gnd), .vdd(vdd), .A(_1084_), .B(_1857_), .Y(_2976_) );
AOI21X1 AOI21X1_258 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(_2959_), .C(_2976_), .Y(_2977_) );
NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(_2968_), .B(_2961_), .Y(_2978_) );
OAI21X1 OAI21X1_1464 ( .gnd(gnd), .vdd(vdd), .A(_2978_), .B(_2958_), .C(_2977_), .Y(_2979_) );
AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(_2979_), .B(_2975_), .Y(_2980_) );
OAI21X1 OAI21X1_1465 ( .gnd(gnd), .vdd(vdd), .A(_2975_), .B(_2979_), .C(digest_valid_new_bF_buf5), .Y(_2981_) );
OAI22X1 OAI22X1_110 ( .gnd(gnd), .vdd(vdd), .A(_1860_), .B(_2006__bF_buf6), .C(_2980_), .D(_2981_), .Y(_3__22_) );
NOR2X1 NOR2X1_572 ( .gnd(gnd), .vdd(vdd), .A(_2973_), .B(_2980_), .Y(_2982_) );
NOR2X1 NOR2X1_573 ( .gnd(gnd), .vdd(vdd), .A(_1205_), .B(_1863_), .Y(_2983_) );
NOR2X1 NOR2X1_574 ( .gnd(gnd), .vdd(vdd), .A(d_reg_23_), .B(_3667__55_), .Y(_2984_) );
NOR2X1 NOR2X1_575 ( .gnd(gnd), .vdd(vdd), .A(_2984_), .B(_2983_), .Y(_2985_) );
XOR2X1 XOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_2982_), .B(_2985_), .Y(_2986_) );
OAI22X1 OAI22X1_111 ( .gnd(gnd), .vdd(vdd), .A(_1863_), .B(_2006__bF_buf5), .C(_2005__bF_buf8), .D(_2986_), .Y(_3__23_) );
NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(_2975_), .B(_2985_), .Y(_2987_) );
NOR2X1 NOR2X1_576 ( .gnd(gnd), .vdd(vdd), .A(_2978_), .B(_2987_), .Y(_2988_) );
NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_2988_), .B(_2955_), .Y(_2989_) );
INVX1 INVX1_979 ( .gnd(gnd), .vdd(vdd), .A(_2989_), .Y(_2990_) );
AOI21X1 AOI21X1_259 ( .gnd(gnd), .vdd(vdd), .A(_2985_), .B(_2973_), .C(_2983_), .Y(_2991_) );
OAI21X1 OAI21X1_1466 ( .gnd(gnd), .vdd(vdd), .A(_2987_), .B(_2977_), .C(_2991_), .Y(_2992_) );
NOR2X1 NOR2X1_577 ( .gnd(gnd), .vdd(vdd), .A(_2992_), .B(_2990_), .Y(_2993_) );
INVX1 INVX1_980 ( .gnd(gnd), .vdd(vdd), .A(_2993_), .Y(_2994_) );
AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(_2957_), .B(_2988_), .Y(_2995_) );
AOI21X1 AOI21X1_260 ( .gnd(gnd), .vdd(vdd), .A(_2923_), .B(_2995_), .C(_2994_), .Y(_2996_) );
NOR2X1 NOR2X1_578 ( .gnd(gnd), .vdd(vdd), .A(_1268_), .B(_1866_), .Y(_2997_) );
NOR2X1 NOR2X1_579 ( .gnd(gnd), .vdd(vdd), .A(d_reg_24_), .B(_3667__56_), .Y(_2998_) );
NOR2X1 NOR2X1_580 ( .gnd(gnd), .vdd(vdd), .A(_2998_), .B(_2997_), .Y(_2999_) );
INVX1 INVX1_981 ( .gnd(gnd), .vdd(vdd), .A(_2999_), .Y(_3000_) );
NOR2X1 NOR2X1_581 ( .gnd(gnd), .vdd(vdd), .A(_3000_), .B(_2996_), .Y(_3001_) );
INVX1 INVX1_982 ( .gnd(gnd), .vdd(vdd), .A(_2996_), .Y(_3002_) );
OAI21X1 OAI21X1_1467 ( .gnd(gnd), .vdd(vdd), .A(_2999_), .B(_3002_), .C(digest_valid_new_bF_buf4), .Y(_3003_) );
OAI22X1 OAI22X1_112 ( .gnd(gnd), .vdd(vdd), .A(_1866_), .B(_2006__bF_buf4), .C(_3001_), .D(_3003_), .Y(_3__24_) );
INVX1 INVX1_983 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .Y(_3004_) );
NOR2X1 NOR2X1_582 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1869_), .Y(_3005_) );
NOR2X1 NOR2X1_583 ( .gnd(gnd), .vdd(vdd), .A(d_reg_25_), .B(_3667__57_), .Y(_3006_) );
OAI21X1 OAI21X1_1468 ( .gnd(gnd), .vdd(vdd), .A(_3005_), .B(_3006_), .C(_3004_), .Y(_3007_) );
NOR2X1 NOR2X1_584 ( .gnd(gnd), .vdd(vdd), .A(_3006_), .B(_3005_), .Y(_3008_) );
OAI21X1 OAI21X1_1469 ( .gnd(gnd), .vdd(vdd), .A(_2997_), .B(_3001_), .C(_3008_), .Y(_3009_) );
OAI21X1 OAI21X1_1470 ( .gnd(gnd), .vdd(vdd), .A(_3001_), .B(_3007_), .C(_3009_), .Y(_3010_) );
OAI22X1 OAI22X1_113 ( .gnd(gnd), .vdd(vdd), .A(_1869_), .B(_2006__bF_buf3), .C(_2005__bF_buf7), .D(_3010_), .Y(_3__25_) );
INVX1 INVX1_984 ( .gnd(gnd), .vdd(vdd), .A(_3008_), .Y(_3011_) );
NOR2X1 NOR2X1_585 ( .gnd(gnd), .vdd(vdd), .A(_3000_), .B(_3011_), .Y(_3012_) );
INVX1 INVX1_985 ( .gnd(gnd), .vdd(vdd), .A(_3012_), .Y(_3013_) );
NOR2X1 NOR2X1_586 ( .gnd(gnd), .vdd(vdd), .A(_3004_), .B(_3011_), .Y(_3014_) );
INVX1 INVX1_986 ( .gnd(gnd), .vdd(vdd), .A(_3014_), .Y(_3015_) );
OAI21X1 OAI21X1_1471 ( .gnd(gnd), .vdd(vdd), .A(_1309_), .B(_1869_), .C(_3015_), .Y(_3016_) );
INVX1 INVX1_987 ( .gnd(gnd), .vdd(vdd), .A(_3016_), .Y(_3017_) );
OAI21X1 OAI21X1_1472 ( .gnd(gnd), .vdd(vdd), .A(_3013_), .B(_2996_), .C(_3017_), .Y(_3018_) );
NOR2X1 NOR2X1_587 ( .gnd(gnd), .vdd(vdd), .A(_1348_), .B(_1872_), .Y(_3019_) );
NOR2X1 NOR2X1_588 ( .gnd(gnd), .vdd(vdd), .A(d_reg_26_), .B(_3667__58_), .Y(_3020_) );
NOR2X1 NOR2X1_589 ( .gnd(gnd), .vdd(vdd), .A(_3020_), .B(_3019_), .Y(_3021_) );
AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(_3018_), .B(_3021_), .Y(_3022_) );
OAI21X1 OAI21X1_1473 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_3018_), .C(digest_valid_new_bF_buf3), .Y(_3023_) );
OAI22X1 OAI22X1_114 ( .gnd(gnd), .vdd(vdd), .A(_1872_), .B(_2006__bF_buf2), .C(_3022_), .D(_3023_), .Y(_3__26_) );
NOR2X1 NOR2X1_590 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(_1876_), .Y(_3024_) );
NOR2X1 NOR2X1_591 ( .gnd(gnd), .vdd(vdd), .A(d_reg_27_), .B(_3667__59_), .Y(_3025_) );
NOR2X1 NOR2X1_592 ( .gnd(gnd), .vdd(vdd), .A(_3025_), .B(_3024_), .Y(_3026_) );
OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(_3022_), .B(_3019_), .Y(_3027_) );
NOR2X1 NOR2X1_593 ( .gnd(gnd), .vdd(vdd), .A(_3026_), .B(_3027_), .Y(_3028_) );
OAI21X1 OAI21X1_1474 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3022_), .C(_3026_), .Y(_3029_) );
NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf2), .B(_3029_), .Y(_3030_) );
OAI22X1 OAI22X1_115 ( .gnd(gnd), .vdd(vdd), .A(_1876_), .B(_2006__bF_buf1), .C(_3030_), .D(_3028_), .Y(_3__27_) );
NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_3021_), .B(_3026_), .Y(_3031_) );
INVX1 INVX1_988 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .Y(_3032_) );
NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_3019_), .B(_3026_), .Y(_3033_) );
OAI21X1 OAI21X1_1475 ( .gnd(gnd), .vdd(vdd), .A(_1875_), .B(_1876_), .C(_3033_), .Y(_3034_) );
AOI21X1 AOI21X1_261 ( .gnd(gnd), .vdd(vdd), .A(_3016_), .B(_3032_), .C(_3034_), .Y(_3035_) );
NOR2X1 NOR2X1_594 ( .gnd(gnd), .vdd(vdd), .A(_3031_), .B(_3013_), .Y(_3036_) );
INVX1 INVX1_989 ( .gnd(gnd), .vdd(vdd), .A(_3036_), .Y(_3037_) );
OAI21X1 OAI21X1_1476 ( .gnd(gnd), .vdd(vdd), .A(_3037_), .B(_2996_), .C(_3035_), .Y(_3038_) );
NOR2X1 NOR2X1_595 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1879_), .Y(_3039_) );
NOR2X1 NOR2X1_596 ( .gnd(gnd), .vdd(vdd), .A(d_reg_28_), .B(_3667__60_), .Y(_3040_) );
NOR2X1 NOR2X1_597 ( .gnd(gnd), .vdd(vdd), .A(_3040_), .B(_3039_), .Y(_3041_) );
NOR2X1 NOR2X1_598 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_3038_), .Y(_3042_) );
NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_3038_), .Y(_3043_) );
NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf1), .B(_3043_), .Y(_3044_) );
OAI21X1 OAI21X1_1477 ( .gnd(gnd), .vdd(vdd), .A(_3667__60_), .B(_3432__bF_buf9), .C(_2005__bF_buf6), .Y(_3045_) );
OAI21X1 OAI21X1_1478 ( .gnd(gnd), .vdd(vdd), .A(_3042_), .B(_3044_), .C(_3045_), .Y(_3__28_) );
OAI21X1 OAI21X1_1479 ( .gnd(gnd), .vdd(vdd), .A(_1436_), .B(_1879_), .C(_3043_), .Y(_3046_) );
NOR2X1 NOR2X1_599 ( .gnd(gnd), .vdd(vdd), .A(_1474_), .B(_1882_), .Y(_3047_) );
NOR2X1 NOR2X1_600 ( .gnd(gnd), .vdd(vdd), .A(d_reg_29_), .B(_3667__61_), .Y(_3048_) );
NOR2X1 NOR2X1_601 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .B(_3047_), .Y(_3049_) );
XNOR2X1 XNOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(_3046_), .B(_3049_), .Y(_3050_) );
OAI22X1 OAI22X1_116 ( .gnd(gnd), .vdd(vdd), .A(_1882_), .B(_2006__bF_buf0), .C(_2005__bF_buf5), .D(_3050_), .Y(_3__29_) );
NOR2X1 NOR2X1_602 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_1885_), .Y(_3051_) );
INVX1 INVX1_990 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .Y(_3052_) );
NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_1526_), .B(_1885_), .Y(_3053_) );
AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(_3052_), .B(_3053_), .Y(_3054_) );
INVX1 INVX1_991 ( .gnd(gnd), .vdd(vdd), .A(_3054_), .Y(_3055_) );
INVX1 INVX1_992 ( .gnd(gnd), .vdd(vdd), .A(_3048_), .Y(_3056_) );
AOI21X1 AOI21X1_262 ( .gnd(gnd), .vdd(vdd), .A(_3039_), .B(_3056_), .C(_3047_), .Y(_3057_) );
INVX1 INVX1_993 ( .gnd(gnd), .vdd(vdd), .A(_3057_), .Y(_3058_) );
AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(_3041_), .B(_3049_), .Y(_3059_) );
AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(_3038_), .B(_3059_), .Y(_3060_) );
NOR2X1 NOR2X1_603 ( .gnd(gnd), .vdd(vdd), .A(_3058_), .B(_3060_), .Y(_3061_) );
AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(_3061_), .B(_3055_), .Y(_3062_) );
OAI21X1 OAI21X1_1480 ( .gnd(gnd), .vdd(vdd), .A(_3055_), .B(_3061_), .C(digest_valid_new_bF_buf0), .Y(_3063_) );
OAI22X1 OAI22X1_117 ( .gnd(gnd), .vdd(vdd), .A(_1885_), .B(_2006__bF_buf8), .C(_3062_), .D(_3063_), .Y(_3__30_) );
INVX1 INVX1_994 ( .gnd(gnd), .vdd(vdd), .A(_3667__63_), .Y(_3064_) );
NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_3059_), .B(_3038_), .Y(_3065_) );
AOI21X1 AOI21X1_263 ( .gnd(gnd), .vdd(vdd), .A(_3065_), .B(_3057_), .C(_3055_), .Y(_3066_) );
XOR2X1 XOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(d_reg_31_), .B(_3667__63_), .Y(_3067_) );
OAI21X1 OAI21X1_1481 ( .gnd(gnd), .vdd(vdd), .A(_3051_), .B(_3066_), .C(_3067_), .Y(_3068_) );
OAI21X1 OAI21X1_1482 ( .gnd(gnd), .vdd(vdd), .A(_3058_), .B(_3060_), .C(_3054_), .Y(_3069_) );
INVX1 INVX1_995 ( .gnd(gnd), .vdd(vdd), .A(_3067_), .Y(_3070_) );
NAND3X1 NAND3X1_306 ( .gnd(gnd), .vdd(vdd), .A(_3052_), .B(_3070_), .C(_3069_), .Y(_3071_) );
NAND3X1 NAND3X1_307 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf8), .B(_3068_), .C(_3071_), .Y(_3072_) );
OAI21X1 OAI21X1_1483 ( .gnd(gnd), .vdd(vdd), .A(_3064_), .B(_2006__bF_buf7), .C(_3072_), .Y(_3__31_) );
XNOR2X1 XNOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(e_reg_0_), .B(_3667__0_), .Y(_3073_) );
OAI22X1 OAI22X1_118 ( .gnd(gnd), .vdd(vdd), .A(_1893_), .B(_2006__bF_buf6), .C(_2005__bF_buf4), .D(_3073_), .Y(_4__0_) );
NOR2X1 NOR2X1_604 ( .gnd(gnd), .vdd(vdd), .A(_1892_), .B(_1893_), .Y(_3074_) );
XOR2X1 XOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(e_reg_1_), .B(_3667__1_), .Y(_3075_) );
XNOR2X1 XNOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(_3075_), .B(_3074_), .Y(_3076_) );
OAI22X1 OAI22X1_119 ( .gnd(gnd), .vdd(vdd), .A(_1897_), .B(_2006__bF_buf5), .C(_2005__bF_buf3), .D(_3076_), .Y(_4__1_) );
NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_3074_), .B(_3075_), .Y(_3077_) );
OAI21X1 OAI21X1_1484 ( .gnd(gnd), .vdd(vdd), .A(_1896_), .B(_1897_), .C(_3077_), .Y(_3078_) );
NOR2X1 NOR2X1_605 ( .gnd(gnd), .vdd(vdd), .A(_1900_), .B(_1901_), .Y(_3079_) );
NOR2X1 NOR2X1_606 ( .gnd(gnd), .vdd(vdd), .A(e_reg_2_), .B(_3667__2_), .Y(_3080_) );
NOR2X1 NOR2X1_607 ( .gnd(gnd), .vdd(vdd), .A(_3080_), .B(_3079_), .Y(_3081_) );
XNOR2X1 XNOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(_3078_), .B(_3081_), .Y(_3082_) );
OAI22X1 OAI22X1_120 ( .gnd(gnd), .vdd(vdd), .A(_1901_), .B(_2006__bF_buf4), .C(_2005__bF_buf2), .D(_3082_), .Y(_4__2_) );
AOI21X1 AOI21X1_264 ( .gnd(gnd), .vdd(vdd), .A(_3078_), .B(_3081_), .C(_3079_), .Y(_3083_) );
NOR2X1 NOR2X1_608 ( .gnd(gnd), .vdd(vdd), .A(_1904_), .B(_1905_), .Y(_3084_) );
NOR2X1 NOR2X1_609 ( .gnd(gnd), .vdd(vdd), .A(e_reg_3_), .B(_3667__3_), .Y(_3085_) );
NOR2X1 NOR2X1_610 ( .gnd(gnd), .vdd(vdd), .A(_3085_), .B(_3084_), .Y(_3086_) );
XOR2X1 XOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_3083_), .B(_3086_), .Y(_3087_) );
OAI22X1 OAI22X1_121 ( .gnd(gnd), .vdd(vdd), .A(_1905_), .B(_2006__bF_buf3), .C(_2005__bF_buf1), .D(_3087_), .Y(_4__3_) );
NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(e_reg_4_), .B(_3667__4_), .Y(_3088_) );
NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(_1909_), .Y(_3089_) );
NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_3089_), .Y(_3090_) );
INVX1 INVX1_996 ( .gnd(gnd), .vdd(vdd), .A(_3090_), .Y(_3091_) );
INVX1 INVX1_997 ( .gnd(gnd), .vdd(vdd), .A(_3084_), .Y(_3092_) );
OAI21X1 OAI21X1_1485 ( .gnd(gnd), .vdd(vdd), .A(_3085_), .B(_3083_), .C(_3092_), .Y(_3093_) );
NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(_3091_), .B(_3093_), .Y(_3094_) );
INVX1 INVX1_998 ( .gnd(gnd), .vdd(vdd), .A(_3093_), .Y(_3095_) );
NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_3090_), .B(_3095_), .Y(_3096_) );
NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3094_), .B(_3096_), .Y(_3097_) );
NOR2X1 NOR2X1_611 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf7), .B(_1910_), .Y(_3098_) );
AOI21X1 AOI21X1_265 ( .gnd(gnd), .vdd(vdd), .A(_3097_), .B(digest_valid_new_bF_buf6), .C(_3098_), .Y(_4__4_) );
OAI21X1 OAI21X1_1486 ( .gnd(gnd), .vdd(vdd), .A(_1908_), .B(_1909_), .C(_3094_), .Y(_3099_) );
NOR2X1 NOR2X1_612 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_1912_), .Y(_3100_) );
NOR2X1 NOR2X1_613 ( .gnd(gnd), .vdd(vdd), .A(e_reg_5_), .B(_3667__5_), .Y(_3101_) );
OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(_3100_), .B(_3101_), .Y(_3102_) );
INVX1 INVX1_999 ( .gnd(gnd), .vdd(vdd), .A(_3102_), .Y(_3103_) );
NOR2X1 NOR2X1_614 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .B(_3099_), .Y(_3104_) );
NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_3103_), .B(_3099_), .Y(_3105_) );
NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf5), .B(_3105_), .Y(_3106_) );
OAI21X1 OAI21X1_1487 ( .gnd(gnd), .vdd(vdd), .A(_3667__5_), .B(_3432__bF_buf8), .C(_2005__bF_buf0), .Y(_3107_) );
OAI21X1 OAI21X1_1488 ( .gnd(gnd), .vdd(vdd), .A(_3104_), .B(_3106_), .C(_3107_), .Y(_4__5_) );
OAI21X1 OAI21X1_1489 ( .gnd(gnd), .vdd(vdd), .A(_72_), .B(_1912_), .C(_3105_), .Y(_3108_) );
XNOR2X1 XNOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(e_reg_6_), .B(_3667__6_), .Y(_3109_) );
INVX1 INVX1_1000 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .Y(_3110_) );
NOR2X1 NOR2X1_615 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .B(_3108_), .Y(_3111_) );
NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_3110_), .B(_3108_), .Y(_3112_) );
NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf4), .B(_3112_), .Y(_3113_) );
OAI21X1 OAI21X1_1490 ( .gnd(gnd), .vdd(vdd), .A(_3667__6_), .B(_3432__bF_buf7), .C(_2005__bF_buf11), .Y(_3114_) );
OAI21X1 OAI21X1_1491 ( .gnd(gnd), .vdd(vdd), .A(_3111_), .B(_3113_), .C(_3114_), .Y(_4__6_) );
OAI21X1 OAI21X1_1492 ( .gnd(gnd), .vdd(vdd), .A(_1915_), .B(_1916_), .C(_3112_), .Y(_3115_) );
INVX1 INVX1_1001 ( .gnd(gnd), .vdd(vdd), .A(_3115_), .Y(_3116_) );
NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(e_reg_7_), .B(_3667__7_), .Y(_3117_) );
NOR2X1 NOR2X1_616 ( .gnd(gnd), .vdd(vdd), .A(e_reg_7_), .B(_3667__7_), .Y(_3118_) );
INVX1 INVX1_1002 ( .gnd(gnd), .vdd(vdd), .A(_3118_), .Y(_3119_) );
NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_3117_), .B(_3119_), .Y(_3120_) );
INVX1 INVX1_1003 ( .gnd(gnd), .vdd(vdd), .A(_3120_), .Y(_3121_) );
NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(_3121_), .B(_3116_), .Y(_3122_) );
INVX1 INVX1_1004 ( .gnd(gnd), .vdd(vdd), .A(_3122_), .Y(_3123_) );
NOR2X1 NOR2X1_617 ( .gnd(gnd), .vdd(vdd), .A(_3121_), .B(_3116_), .Y(_3124_) );
OAI21X1 OAI21X1_1493 ( .gnd(gnd), .vdd(vdd), .A(_3124_), .B(_3123_), .C(digest_valid_new_bF_buf3), .Y(_3125_) );
OAI21X1 OAI21X1_1494 ( .gnd(gnd), .vdd(vdd), .A(_3667__7_), .B(_3432__bF_buf6), .C(_2005__bF_buf10), .Y(_3126_) );
NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3126_), .B(_3125_), .Y(_4__7_) );
NOR2X1 NOR2X1_618 ( .gnd(gnd), .vdd(vdd), .A(_1921_), .B(_1922_), .Y(_3127_) );
NOR2X1 NOR2X1_619 ( .gnd(gnd), .vdd(vdd), .A(e_reg_8_), .B(_3667__8_), .Y(_3128_) );
NOR2X1 NOR2X1_620 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_3127_), .Y(_3129_) );
NOR2X1 NOR2X1_621 ( .gnd(gnd), .vdd(vdd), .A(_3088_), .B(_3102_), .Y(_3130_) );
OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(_3130_), .B(_3100_), .Y(_3131_) );
NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(e_reg_6_), .B(_3667__6_), .Y(_3132_) );
OAI21X1 OAI21X1_1495 ( .gnd(gnd), .vdd(vdd), .A(_3132_), .B(_3118_), .C(_3117_), .Y(_3133_) );
NOR2X1 NOR2X1_622 ( .gnd(gnd), .vdd(vdd), .A(_3109_), .B(_3120_), .Y(_3134_) );
AOI21X1 AOI21X1_266 ( .gnd(gnd), .vdd(vdd), .A(_3134_), .B(_3131_), .C(_3133_), .Y(_3135_) );
NAND3X1 NAND3X1_308 ( .gnd(gnd), .vdd(vdd), .A(_3091_), .B(_3134_), .C(_3103_), .Y(_3136_) );
OAI21X1 OAI21X1_1496 ( .gnd(gnd), .vdd(vdd), .A(_3136_), .B(_3095_), .C(_3135_), .Y(_3137_) );
NOR2X1 NOR2X1_623 ( .gnd(gnd), .vdd(vdd), .A(_3129_), .B(_3137_), .Y(_3138_) );
INVX1 INVX1_1005 ( .gnd(gnd), .vdd(vdd), .A(_3129_), .Y(_3139_) );
INVX1 INVX1_1006 ( .gnd(gnd), .vdd(vdd), .A(_3137_), .Y(_3140_) );
OAI21X1 OAI21X1_1497 ( .gnd(gnd), .vdd(vdd), .A(_3139_), .B(_3140_), .C(digest_valid_new_bF_buf2), .Y(_3141_) );
OAI21X1 OAI21X1_1498 ( .gnd(gnd), .vdd(vdd), .A(_3667__8_), .B(_3432__bF_buf5), .C(_2005__bF_buf9), .Y(_3142_) );
OAI21X1 OAI21X1_1499 ( .gnd(gnd), .vdd(vdd), .A(_3138_), .B(_3141_), .C(_3142_), .Y(_4__8_) );
NOR2X1 NOR2X1_624 ( .gnd(gnd), .vdd(vdd), .A(_1925_), .B(_1926_), .Y(_3143_) );
NOR2X1 NOR2X1_625 ( .gnd(gnd), .vdd(vdd), .A(e_reg_9_), .B(_3667__9_), .Y(_3144_) );
OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .B(_3144_), .Y(_3145_) );
INVX1 INVX1_1007 ( .gnd(gnd), .vdd(vdd), .A(_3145_), .Y(_3146_) );
INVX1 INVX1_1008 ( .gnd(gnd), .vdd(vdd), .A(_3127_), .Y(_3147_) );
OAI21X1 OAI21X1_1500 ( .gnd(gnd), .vdd(vdd), .A(_3128_), .B(_3140_), .C(_3147_), .Y(_3148_) );
NOR2X1 NOR2X1_626 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(_3148_), .Y(_3149_) );
NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(_3146_), .B(_3148_), .Y(_3150_) );
NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf1), .B(_3150_), .Y(_3151_) );
OAI22X1 OAI22X1_122 ( .gnd(gnd), .vdd(vdd), .A(_1926_), .B(_2006__bF_buf2), .C(_3149_), .D(_3151_), .Y(_4__9_) );
INVX1 INVX1_1009 ( .gnd(gnd), .vdd(vdd), .A(_3143_), .Y(_3152_) );
NOR2X1 NOR2X1_627 ( .gnd(gnd), .vdd(vdd), .A(_1929_), .B(_1930_), .Y(_3153_) );
NOR2X1 NOR2X1_628 ( .gnd(gnd), .vdd(vdd), .A(e_reg_10_), .B(_3667__10_), .Y(_3154_) );
OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(_3153_), .B(_3154_), .Y(_3155_) );
AOI21X1 AOI21X1_267 ( .gnd(gnd), .vdd(vdd), .A(_3150_), .B(_3152_), .C(_3155_), .Y(_3156_) );
OAI21X1 OAI21X1_1501 ( .gnd(gnd), .vdd(vdd), .A(_1925_), .B(_1926_), .C(_3150_), .Y(_3157_) );
INVX1 INVX1_1010 ( .gnd(gnd), .vdd(vdd), .A(_3155_), .Y(_3158_) );
OAI21X1 OAI21X1_1502 ( .gnd(gnd), .vdd(vdd), .A(_3158_), .B(_3157_), .C(digest_valid_new_bF_buf0), .Y(_3159_) );
OAI22X1 OAI22X1_123 ( .gnd(gnd), .vdd(vdd), .A(_1930_), .B(_2006__bF_buf1), .C(_3156_), .D(_3159_), .Y(_4__10_) );
NOR2X1 NOR2X1_629 ( .gnd(gnd), .vdd(vdd), .A(_3153_), .B(_3156_), .Y(_3160_) );
XOR2X1 XOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(e_reg_11_), .B(_3667__11_), .Y(_3161_) );
INVX1 INVX1_1011 ( .gnd(gnd), .vdd(vdd), .A(_3161_), .Y(_3162_) );
XNOR2X1 XNOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(_3160_), .B(_3162_), .Y(_3163_) );
OAI22X1 OAI22X1_124 ( .gnd(gnd), .vdd(vdd), .A(_1934_), .B(_2006__bF_buf0), .C(_2005__bF_buf8), .D(_3163_), .Y(_4__11_) );
OAI21X1 OAI21X1_1503 ( .gnd(gnd), .vdd(vdd), .A(_3144_), .B(_3147_), .C(_3152_), .Y(_3164_) );
NOR2X1 NOR2X1_630 ( .gnd(gnd), .vdd(vdd), .A(_3162_), .B(_3155_), .Y(_3165_) );
OAI21X1 OAI21X1_1504 ( .gnd(gnd), .vdd(vdd), .A(e_reg_11_), .B(_3667__11_), .C(_3153_), .Y(_3166_) );
OAI21X1 OAI21X1_1505 ( .gnd(gnd), .vdd(vdd), .A(_1933_), .B(_1934_), .C(_3166_), .Y(_3167_) );
AOI21X1 AOI21X1_268 ( .gnd(gnd), .vdd(vdd), .A(_3165_), .B(_3164_), .C(_3167_), .Y(_3168_) );
NAND3X1 NAND3X1_309 ( .gnd(gnd), .vdd(vdd), .A(_3129_), .B(_3146_), .C(_3165_), .Y(_3169_) );
OAI21X1 OAI21X1_1506 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .B(_3140_), .C(_3168_), .Y(_3170_) );
NOR2X1 NOR2X1_631 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .B(_1938_), .Y(_3171_) );
NOR2X1 NOR2X1_632 ( .gnd(gnd), .vdd(vdd), .A(e_reg_12_), .B(_3667__12_), .Y(_3172_) );
NOR2X1 NOR2X1_633 ( .gnd(gnd), .vdd(vdd), .A(_3172_), .B(_3171_), .Y(_3173_) );
NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_3173_), .B(_3170_), .Y(_3174_) );
INVX1 INVX1_1012 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .Y(_3175_) );
OAI21X1 OAI21X1_1507 ( .gnd(gnd), .vdd(vdd), .A(_3173_), .B(_3170_), .C(digest_valid_new_bF_buf8), .Y(_3176_) );
OAI22X1 OAI22X1_125 ( .gnd(gnd), .vdd(vdd), .A(_1938_), .B(_2006__bF_buf8), .C(_3176_), .D(_3175_), .Y(_4__12_) );
OAI21X1 OAI21X1_1508 ( .gnd(gnd), .vdd(vdd), .A(_1937_), .B(_1938_), .C(_3174_), .Y(_3177_) );
NOR2X1 NOR2X1_634 ( .gnd(gnd), .vdd(vdd), .A(_1941_), .B(_1942_), .Y(_3178_) );
NOR2X1 NOR2X1_635 ( .gnd(gnd), .vdd(vdd), .A(e_reg_13_), .B(_3667__13_), .Y(_3179_) );
NOR2X1 NOR2X1_636 ( .gnd(gnd), .vdd(vdd), .A(_3179_), .B(_3178_), .Y(_3180_) );
XNOR2X1 XNOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(_3177_), .B(_3180_), .Y(_3181_) );
OAI21X1 OAI21X1_1509 ( .gnd(gnd), .vdd(vdd), .A(_3667__13_), .B(_3432__bF_buf4), .C(_2005__bF_buf7), .Y(_3182_) );
OAI21X1 OAI21X1_1510 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf6), .B(_3181_), .C(_3182_), .Y(_4__13_) );
NOR2X1 NOR2X1_637 ( .gnd(gnd), .vdd(vdd), .A(_1945_), .B(_1946_), .Y(_3183_) );
NOR2X1 NOR2X1_638 ( .gnd(gnd), .vdd(vdd), .A(e_reg_14_), .B(_3667__14_), .Y(_3184_) );
NOR2X1 NOR2X1_639 ( .gnd(gnd), .vdd(vdd), .A(_3184_), .B(_3183_), .Y(_3185_) );
NOR2X1 NOR2X1_640 ( .gnd(gnd), .vdd(vdd), .A(_3171_), .B(_3178_), .Y(_3186_) );
AOI21X1 AOI21X1_269 ( .gnd(gnd), .vdd(vdd), .A(_3174_), .B(_3186_), .C(_3179_), .Y(_3187_) );
NOR2X1 NOR2X1_641 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .B(_3187_), .Y(_3188_) );
INVX1 INVX1_1013 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .Y(_3189_) );
INVX1 INVX1_1014 ( .gnd(gnd), .vdd(vdd), .A(_3187_), .Y(_3190_) );
OAI21X1 OAI21X1_1511 ( .gnd(gnd), .vdd(vdd), .A(_3189_), .B(_3190_), .C(digest_valid_new_bF_buf7), .Y(_3191_) );
OAI21X1 OAI21X1_1512 ( .gnd(gnd), .vdd(vdd), .A(_3667__14_), .B(_3432__bF_buf3), .C(_2005__bF_buf5), .Y(_3192_) );
OAI21X1 OAI21X1_1513 ( .gnd(gnd), .vdd(vdd), .A(_3188_), .B(_3191_), .C(_3192_), .Y(_4__14_) );
AOI21X1 AOI21X1_270 ( .gnd(gnd), .vdd(vdd), .A(_3187_), .B(_3185_), .C(_3183_), .Y(_3193_) );
NOR2X1 NOR2X1_642 ( .gnd(gnd), .vdd(vdd), .A(_1949_), .B(_1950_), .Y(_3194_) );
NOR2X1 NOR2X1_643 ( .gnd(gnd), .vdd(vdd), .A(e_reg_15_), .B(_3667__15_), .Y(_3195_) );
NOR2X1 NOR2X1_644 ( .gnd(gnd), .vdd(vdd), .A(_3195_), .B(_3194_), .Y(_3196_) );
XOR2X1 XOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_3193_), .B(_3196_), .Y(_3197_) );
OAI21X1 OAI21X1_1514 ( .gnd(gnd), .vdd(vdd), .A(_3667__15_), .B(_3432__bF_buf2), .C(_2005__bF_buf4), .Y(_3198_) );
OAI21X1 OAI21X1_1515 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf3), .B(_3197_), .C(_3198_), .Y(_4__15_) );
NOR2X1 NOR2X1_645 ( .gnd(gnd), .vdd(vdd), .A(_807_), .B(_1953_), .Y(_3199_) );
NOR2X1 NOR2X1_646 ( .gnd(gnd), .vdd(vdd), .A(e_reg_16_), .B(_3667__16_), .Y(_3200_) );
NOR2X1 NOR2X1_647 ( .gnd(gnd), .vdd(vdd), .A(_3200_), .B(_3199_), .Y(_3201_) );
AOI21X1 AOI21X1_271 ( .gnd(gnd), .vdd(vdd), .A(_3180_), .B(_3171_), .C(_3178_), .Y(_3202_) );
NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_3185_), .B(_3196_), .Y(_3203_) );
AOI21X1 AOI21X1_272 ( .gnd(gnd), .vdd(vdd), .A(_3196_), .B(_3183_), .C(_3194_), .Y(_3204_) );
OAI21X1 OAI21X1_1516 ( .gnd(gnd), .vdd(vdd), .A(_3203_), .B(_3202_), .C(_3204_), .Y(_3205_) );
INVX1 INVX1_1015 ( .gnd(gnd), .vdd(vdd), .A(_3205_), .Y(_3206_) );
NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_3173_), .B(_3180_), .Y(_3207_) );
NOR2X1 NOR2X1_648 ( .gnd(gnd), .vdd(vdd), .A(_3207_), .B(_3203_), .Y(_3208_) );
INVX1 INVX1_1016 ( .gnd(gnd), .vdd(vdd), .A(_3208_), .Y(_3209_) );
OAI21X1 OAI21X1_1517 ( .gnd(gnd), .vdd(vdd), .A(_3209_), .B(_3168_), .C(_3206_), .Y(_3210_) );
NOR2X1 NOR2X1_649 ( .gnd(gnd), .vdd(vdd), .A(_3169_), .B(_3209_), .Y(_3211_) );
AOI21X1 AOI21X1_273 ( .gnd(gnd), .vdd(vdd), .A(_3137_), .B(_3211_), .C(_3210_), .Y(_3212_) );
INVX1 INVX1_1017 ( .gnd(gnd), .vdd(vdd), .A(_3212_), .Y(_3213_) );
NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_3201_), .B(_3213_), .Y(_3214_) );
INVX1 INVX1_1018 ( .gnd(gnd), .vdd(vdd), .A(_3214_), .Y(_3215_) );
OAI21X1 OAI21X1_1518 ( .gnd(gnd), .vdd(vdd), .A(_3201_), .B(_3213_), .C(digest_valid_new_bF_buf6), .Y(_3216_) );
OAI22X1 OAI22X1_126 ( .gnd(gnd), .vdd(vdd), .A(_1953_), .B(_2006__bF_buf7), .C(_3216_), .D(_3215_), .Y(_4__16_) );
INVX1 INVX1_1019 ( .gnd(gnd), .vdd(vdd), .A(_3199_), .Y(_3217_) );
OAI21X1 OAI21X1_1519 ( .gnd(gnd), .vdd(vdd), .A(_3200_), .B(_3212_), .C(_3217_), .Y(_3218_) );
NOR2X1 NOR2X1_650 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_1957_), .Y(_3219_) );
NOR2X1 NOR2X1_651 ( .gnd(gnd), .vdd(vdd), .A(e_reg_17_), .B(_3667__17_), .Y(_3220_) );
NOR2X1 NOR2X1_652 ( .gnd(gnd), .vdd(vdd), .A(_3220_), .B(_3219_), .Y(_3221_) );
XNOR2X1 XNOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(_3218_), .B(_3221_), .Y(_3222_) );
OAI21X1 OAI21X1_1520 ( .gnd(gnd), .vdd(vdd), .A(_3667__17_), .B(_3432__bF_buf1), .C(_2005__bF_buf2), .Y(_3223_) );
OAI21X1 OAI21X1_1521 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf1), .B(_3222_), .C(_3223_), .Y(_4__17_) );
NOR2X1 NOR2X1_653 ( .gnd(gnd), .vdd(vdd), .A(_919_), .B(_1960_), .Y(_3224_) );
NOR2X1 NOR2X1_654 ( .gnd(gnd), .vdd(vdd), .A(e_reg_18_), .B(_3667__18_), .Y(_3225_) );
NOR2X1 NOR2X1_655 ( .gnd(gnd), .vdd(vdd), .A(_3225_), .B(_3224_), .Y(_3226_) );
INVX1 INVX1_1020 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .Y(_3227_) );
INVX1 INVX1_1021 ( .gnd(gnd), .vdd(vdd), .A(_3220_), .Y(_3228_) );
OAI21X1 OAI21X1_1522 ( .gnd(gnd), .vdd(vdd), .A(_1956_), .B(_1957_), .C(_3217_), .Y(_3229_) );
OAI21X1 OAI21X1_1523 ( .gnd(gnd), .vdd(vdd), .A(_3229_), .B(_3215_), .C(_3228_), .Y(_3230_) );
NOR2X1 NOR2X1_656 ( .gnd(gnd), .vdd(vdd), .A(_3227_), .B(_3230_), .Y(_3231_) );
OAI21X1 OAI21X1_1524 ( .gnd(gnd), .vdd(vdd), .A(e_reg_17_), .B(_3667__17_), .C(_3229_), .Y(_3232_) );
NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_3201_), .B(_3221_), .Y(_3233_) );
OAI21X1 OAI21X1_1525 ( .gnd(gnd), .vdd(vdd), .A(_3233_), .B(_3212_), .C(_3232_), .Y(_3234_) );
OAI21X1 OAI21X1_1526 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_3234_), .C(digest_valid_new_bF_buf5), .Y(_3235_) );
OAI22X1 OAI22X1_127 ( .gnd(gnd), .vdd(vdd), .A(_1960_), .B(_2006__bF_buf6), .C(_3235_), .D(_3231_), .Y(_4__18_) );
NOR2X1 NOR2X1_657 ( .gnd(gnd), .vdd(vdd), .A(_1963_), .B(_1964_), .Y(_3236_) );
NOR2X1 NOR2X1_658 ( .gnd(gnd), .vdd(vdd), .A(e_reg_19_), .B(_3667__19_), .Y(_3237_) );
NOR2X1 NOR2X1_659 ( .gnd(gnd), .vdd(vdd), .A(_3237_), .B(_3236_), .Y(_3238_) );
OAI21X1 OAI21X1_1527 ( .gnd(gnd), .vdd(vdd), .A(_3224_), .B(_3231_), .C(_3238_), .Y(_3239_) );
NOR2X1 NOR2X1_660 ( .gnd(gnd), .vdd(vdd), .A(_3224_), .B(_3231_), .Y(_3240_) );
OAI21X1 OAI21X1_1528 ( .gnd(gnd), .vdd(vdd), .A(_3236_), .B(_3237_), .C(_3240_), .Y(_3241_) );
NAND3X1 NAND3X1_310 ( .gnd(gnd), .vdd(vdd), .A(digest_valid_new_bF_buf4), .B(_3239_), .C(_3241_), .Y(_3242_) );
OAI21X1 OAI21X1_1529 ( .gnd(gnd), .vdd(vdd), .A(_1964_), .B(_2006__bF_buf5), .C(_3242_), .Y(_4__19_) );
NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(_3226_), .B(_3238_), .Y(_3243_) );
AOI21X1 AOI21X1_274 ( .gnd(gnd), .vdd(vdd), .A(_3238_), .B(_3224_), .C(_3236_), .Y(_3244_) );
OAI21X1 OAI21X1_1530 ( .gnd(gnd), .vdd(vdd), .A(_3243_), .B(_3232_), .C(_3244_), .Y(_3245_) );
NOR2X1 NOR2X1_661 ( .gnd(gnd), .vdd(vdd), .A(_3233_), .B(_3243_), .Y(_3246_) );
AOI21X1 AOI21X1_275 ( .gnd(gnd), .vdd(vdd), .A(_3213_), .B(_3246_), .C(_3245_), .Y(_3247_) );
NOR2X1 NOR2X1_662 ( .gnd(gnd), .vdd(vdd), .A(_1967_), .B(_1968_), .Y(_3248_) );
NOR2X1 NOR2X1_663 ( .gnd(gnd), .vdd(vdd), .A(e_reg_20_), .B(_3667__20_), .Y(_3249_) );
NOR2X1 NOR2X1_664 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .B(_3248_), .Y(_3250_) );
XOR2X1 XOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(_3247_), .B(_3250_), .Y(_3251_) );
OAI21X1 OAI21X1_1531 ( .gnd(gnd), .vdd(vdd), .A(_3667__20_), .B(_3432__bF_buf0), .C(_2005__bF_buf0), .Y(_3252_) );
OAI21X1 OAI21X1_1532 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf11), .B(_3251_), .C(_3252_), .Y(_4__20_) );
NOR2X1 NOR2X1_665 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1972_), .Y(_3253_) );
NOR2X1 NOR2X1_666 ( .gnd(gnd), .vdd(vdd), .A(e_reg_21_), .B(_3667__21_), .Y(_3254_) );
NOR2X1 NOR2X1_667 ( .gnd(gnd), .vdd(vdd), .A(_3254_), .B(_3253_), .Y(_3255_) );
INVX1 INVX1_1022 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .Y(_3256_) );
OAI21X1 OAI21X1_1533 ( .gnd(gnd), .vdd(vdd), .A(_3249_), .B(_3247_), .C(_3256_), .Y(_3257_) );
NOR2X1 NOR2X1_668 ( .gnd(gnd), .vdd(vdd), .A(_3255_), .B(_3257_), .Y(_3258_) );
NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_3250_), .B(_3255_), .Y(_3259_) );
NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_3248_), .B(_3255_), .Y(_3260_) );
INVX1 INVX1_1023 ( .gnd(gnd), .vdd(vdd), .A(_3260_), .Y(_3261_) );
NOR2X1 NOR2X1_669 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf10), .B(_3261_), .Y(_3262_) );
OAI21X1 OAI21X1_1534 ( .gnd(gnd), .vdd(vdd), .A(_3259_), .B(_3247_), .C(_3262_), .Y(_3263_) );
OAI22X1 OAI22X1_128 ( .gnd(gnd), .vdd(vdd), .A(_1972_), .B(_2006__bF_buf4), .C(_3263_), .D(_3258_), .Y(_4__21_) );
NOR2X1 NOR2X1_670 ( .gnd(gnd), .vdd(vdd), .A(_3259_), .B(_3247_), .Y(_3264_) );
OAI21X1 OAI21X1_1535 ( .gnd(gnd), .vdd(vdd), .A(_1971_), .B(_1972_), .C(_3260_), .Y(_3265_) );
NOR2X1 NOR2X1_671 ( .gnd(gnd), .vdd(vdd), .A(_3265_), .B(_3264_), .Y(_3266_) );
INVX1 INVX1_1024 ( .gnd(gnd), .vdd(vdd), .A(_3266_), .Y(_3267_) );
NOR2X1 NOR2X1_672 ( .gnd(gnd), .vdd(vdd), .A(_1157_), .B(_1975_), .Y(_3268_) );
NOR2X1 NOR2X1_673 ( .gnd(gnd), .vdd(vdd), .A(e_reg_22_), .B(_3667__22_), .Y(_3269_) );
NOR2X1 NOR2X1_674 ( .gnd(gnd), .vdd(vdd), .A(_3269_), .B(_3268_), .Y(_3270_) );
NOR2X1 NOR2X1_675 ( .gnd(gnd), .vdd(vdd), .A(_3270_), .B(_3267_), .Y(_3271_) );
INVX1 INVX1_1025 ( .gnd(gnd), .vdd(vdd), .A(_3270_), .Y(_3272_) );
OAI21X1 OAI21X1_1536 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3266_), .C(digest_valid_new_bF_buf3), .Y(_3273_) );
OAI21X1 OAI21X1_1537 ( .gnd(gnd), .vdd(vdd), .A(_3667__22_), .B(_3432__bF_buf11), .C(_2005__bF_buf9), .Y(_3274_) );
OAI21X1 OAI21X1_1538 ( .gnd(gnd), .vdd(vdd), .A(_3273_), .B(_3271_), .C(_3274_), .Y(_4__22_) );
AOI21X1 AOI21X1_276 ( .gnd(gnd), .vdd(vdd), .A(_3267_), .B(_3270_), .C(_3268_), .Y(_3275_) );
NOR2X1 NOR2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_1215_), .B(_1978_), .Y(_3276_) );
NOR2X1 NOR2X1_677 ( .gnd(gnd), .vdd(vdd), .A(e_reg_23_), .B(_3667__23_), .Y(_3277_) );
NOR2X1 NOR2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_3277_), .B(_3276_), .Y(_3278_) );
INVX1 INVX1_1026 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .Y(_3279_) );
XNOR2X1 XNOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(_3275_), .B(_3279_), .Y(_3280_) );
OAI21X1 OAI21X1_1539 ( .gnd(gnd), .vdd(vdd), .A(_3667__23_), .B(_3432__bF_buf10), .C(_2005__bF_buf8), .Y(_3281_) );
OAI21X1 OAI21X1_1540 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf7), .B(_3280_), .C(_3281_), .Y(_4__23_) );
NOR2X1 NOR2X1_679 ( .gnd(gnd), .vdd(vdd), .A(_3272_), .B(_3279_), .Y(_3282_) );
INVX1 INVX1_1027 ( .gnd(gnd), .vdd(vdd), .A(_3282_), .Y(_3283_) );
NOR2X1 NOR2X1_680 ( .gnd(gnd), .vdd(vdd), .A(_3259_), .B(_3283_), .Y(_3284_) );
NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(_3245_), .B(_3284_), .Y(_3285_) );
OAI21X1 OAI21X1_1541 ( .gnd(gnd), .vdd(vdd), .A(_3253_), .B(_3261_), .C(_3282_), .Y(_3286_) );
AOI21X1 AOI21X1_277 ( .gnd(gnd), .vdd(vdd), .A(_3278_), .B(_3268_), .C(_3276_), .Y(_3287_) );
NAND3X1 NAND3X1_311 ( .gnd(gnd), .vdd(vdd), .A(_3286_), .B(_3287_), .C(_3285_), .Y(_3288_) );
NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(_3246_), .B(_3284_), .Y(_3289_) );
NOR2X1 NOR2X1_681 ( .gnd(gnd), .vdd(vdd), .A(_3289_), .B(_3212_), .Y(_3290_) );
NOR2X1 NOR2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_3288_), .B(_3290_), .Y(_3291_) );
INVX1 INVX1_1028 ( .gnd(gnd), .vdd(vdd), .A(_3291_), .Y(_3292_) );
NOR2X1 NOR2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_1280_), .B(_1981_), .Y(_3293_) );
NOR2X1 NOR2X1_684 ( .gnd(gnd), .vdd(vdd), .A(e_reg_24_), .B(_3667__24_), .Y(_3294_) );
NOR2X1 NOR2X1_685 ( .gnd(gnd), .vdd(vdd), .A(_3294_), .B(_3293_), .Y(_3295_) );
NOR2X1 NOR2X1_686 ( .gnd(gnd), .vdd(vdd), .A(_3295_), .B(_3292_), .Y(_3296_) );
INVX1 INVX1_1029 ( .gnd(gnd), .vdd(vdd), .A(_3295_), .Y(_3297_) );
OAI21X1 OAI21X1_1542 ( .gnd(gnd), .vdd(vdd), .A(_3297_), .B(_3291_), .C(digest_valid_new_bF_buf2), .Y(_3298_) );
OAI21X1 OAI21X1_1543 ( .gnd(gnd), .vdd(vdd), .A(_3667__24_), .B(_3432__bF_buf9), .C(_2005__bF_buf6), .Y(_3299_) );
OAI21X1 OAI21X1_1544 ( .gnd(gnd), .vdd(vdd), .A(_3298_), .B(_3296_), .C(_3299_), .Y(_4__24_) );
AOI21X1 AOI21X1_278 ( .gnd(gnd), .vdd(vdd), .A(_3292_), .B(_3295_), .C(_3293_), .Y(_3300_) );
NOR2X1 NOR2X1_687 ( .gnd(gnd), .vdd(vdd), .A(_1359_), .B(_1984_), .Y(_3301_) );
NOR2X1 NOR2X1_688 ( .gnd(gnd), .vdd(vdd), .A(e_reg_25_), .B(_3667__25_), .Y(_3302_) );
NOR2X1 NOR2X1_689 ( .gnd(gnd), .vdd(vdd), .A(_3302_), .B(_3301_), .Y(_3303_) );
INVX1 INVX1_1030 ( .gnd(gnd), .vdd(vdd), .A(_3303_), .Y(_3304_) );
XNOR2X1 XNOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(_3300_), .B(_3304_), .Y(_3305_) );
OAI21X1 OAI21X1_1545 ( .gnd(gnd), .vdd(vdd), .A(_3667__25_), .B(_3432__bF_buf8), .C(_2005__bF_buf5), .Y(_3306_) );
OAI21X1 OAI21X1_1546 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf4), .B(_3305_), .C(_3306_), .Y(_4__25_) );
NOR2X1 NOR2X1_690 ( .gnd(gnd), .vdd(vdd), .A(_3297_), .B(_3304_), .Y(_3307_) );
INVX1 INVX1_1031 ( .gnd(gnd), .vdd(vdd), .A(_3307_), .Y(_3308_) );
AOI21X1 AOI21X1_279 ( .gnd(gnd), .vdd(vdd), .A(_3303_), .B(_3293_), .C(_3301_), .Y(_3309_) );
OAI21X1 OAI21X1_1547 ( .gnd(gnd), .vdd(vdd), .A(_3308_), .B(_3291_), .C(_3309_), .Y(_3310_) );
NOR2X1 NOR2X1_691 ( .gnd(gnd), .vdd(vdd), .A(_1363_), .B(_1987_), .Y(_3311_) );
NOR2X1 NOR2X1_692 ( .gnd(gnd), .vdd(vdd), .A(e_reg_26_), .B(_3667__26_), .Y(_3312_) );
NOR2X1 NOR2X1_693 ( .gnd(gnd), .vdd(vdd), .A(_3312_), .B(_3311_), .Y(_3313_) );
AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(_3310_), .B(_3313_), .Y(_3314_) );
OAI21X1 OAI21X1_1548 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .B(_3310_), .C(digest_valid_new_bF_buf1), .Y(_3315_) );
OAI22X1 OAI22X1_129 ( .gnd(gnd), .vdd(vdd), .A(_1987_), .B(_2006__bF_buf3), .C(_3314_), .D(_3315_), .Y(_4__26_) );
INVX1 INVX1_1032 ( .gnd(gnd), .vdd(vdd), .A(_3311_), .Y(_3316_) );
NOR2X1 NOR2X1_694 ( .gnd(gnd), .vdd(vdd), .A(_1406_), .B(_1990_), .Y(_3317_) );
NOR2X1 NOR2X1_695 ( .gnd(gnd), .vdd(vdd), .A(e_reg_27_), .B(_3667__27_), .Y(_3318_) );
OAI21X1 OAI21X1_1549 ( .gnd(gnd), .vdd(vdd), .A(_3317_), .B(_3318_), .C(_3316_), .Y(_3319_) );
NOR2X1 NOR2X1_696 ( .gnd(gnd), .vdd(vdd), .A(_3318_), .B(_3317_), .Y(_3320_) );
OAI21X1 OAI21X1_1550 ( .gnd(gnd), .vdd(vdd), .A(_3311_), .B(_3314_), .C(_3320_), .Y(_3321_) );
OAI21X1 OAI21X1_1551 ( .gnd(gnd), .vdd(vdd), .A(_3314_), .B(_3319_), .C(_3321_), .Y(_3322_) );
OAI22X1 OAI22X1_130 ( .gnd(gnd), .vdd(vdd), .A(_1990_), .B(_2006__bF_buf2), .C(_2005__bF_buf3), .D(_3322_), .Y(_4__27_) );
AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(_3313_), .B(_3320_), .Y(_3323_) );
AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(_3310_), .B(_3323_), .Y(_3324_) );
AOI21X1 AOI21X1_280 ( .gnd(gnd), .vdd(vdd), .A(_3320_), .B(_3311_), .C(_3317_), .Y(_3325_) );
INVX1 INVX1_1033 ( .gnd(gnd), .vdd(vdd), .A(_3325_), .Y(_3326_) );
NOR2X1 NOR2X1_697 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .B(_1993_), .Y(_3327_) );
NOR2X1 NOR2X1_698 ( .gnd(gnd), .vdd(vdd), .A(e_reg_28_), .B(_3667__28_), .Y(_3328_) );
NOR2X1 NOR2X1_699 ( .gnd(gnd), .vdd(vdd), .A(_3328_), .B(_3327_), .Y(_3329_) );
OAI21X1 OAI21X1_1552 ( .gnd(gnd), .vdd(vdd), .A(_3326_), .B(_3324_), .C(_3329_), .Y(_3330_) );
NOR2X1 NOR2X1_700 ( .gnd(gnd), .vdd(vdd), .A(_3326_), .B(_3324_), .Y(_3331_) );
OAI21X1 OAI21X1_1553 ( .gnd(gnd), .vdd(vdd), .A(_3327_), .B(_3328_), .C(_3331_), .Y(_3332_) );
NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(_3330_), .B(_3332_), .Y(_3333_) );
OAI22X1 OAI22X1_131 ( .gnd(gnd), .vdd(vdd), .A(_1993_), .B(_2006__bF_buf1), .C(_2005__bF_buf2), .D(_3333_), .Y(_4__28_) );
OAI21X1 OAI21X1_1554 ( .gnd(gnd), .vdd(vdd), .A(_1484_), .B(_1993_), .C(_3330_), .Y(_3334_) );
NOR2X1 NOR2X1_701 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_1996_), .Y(_3335_) );
NOR2X1 NOR2X1_702 ( .gnd(gnd), .vdd(vdd), .A(e_reg_29_), .B(_3667__29_), .Y(_3336_) );
NOR2X1 NOR2X1_703 ( .gnd(gnd), .vdd(vdd), .A(_3336_), .B(_3335_), .Y(_3337_) );
XNOR2X1 XNOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(_3334_), .B(_3337_), .Y(_3338_) );
OAI22X1 OAI22X1_132 ( .gnd(gnd), .vdd(vdd), .A(_1996_), .B(_2006__bF_buf0), .C(_2005__bF_buf1), .D(_3338_), .Y(_4__29_) );
NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(e_reg_30_), .B(_3667__30_), .Y(_3339_) );
OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(e_reg_30_), .B(_3667__30_), .Y(_3340_) );
AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(_3340_), .B(_3339_), .Y(_3341_) );
OAI21X1 OAI21X1_1555 ( .gnd(gnd), .vdd(vdd), .A(e_reg_29_), .B(_3667__29_), .C(_3334_), .Y(_3342_) );
OAI21X1 OAI21X1_1556 ( .gnd(gnd), .vdd(vdd), .A(_1488_), .B(_1996_), .C(_3342_), .Y(_3343_) );
XNOR2X1 XNOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(_3343_), .B(_3341_), .Y(_3344_) );
OAI21X1 OAI21X1_1557 ( .gnd(gnd), .vdd(vdd), .A(_3667__30_), .B(_3432__bF_buf7), .C(_2005__bF_buf0), .Y(_3345_) );
OAI21X1 OAI21X1_1558 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf11), .B(_3344_), .C(_3345_), .Y(_4__30_) );
NOR2X1 NOR2X1_704 ( .gnd(gnd), .vdd(vdd), .A(_3667__31_), .B(_3432__bF_buf6), .Y(_3346_) );
INVX1 INVX1_1034 ( .gnd(gnd), .vdd(vdd), .A(_3339_), .Y(_3347_) );
AOI21X1 AOI21X1_281 ( .gnd(gnd), .vdd(vdd), .A(_3343_), .B(_3341_), .C(_3347_), .Y(_3348_) );
XNOR2X1 XNOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(e_reg_31_), .B(_3667__31_), .Y(_3349_) );
INVX1 INVX1_1035 ( .gnd(gnd), .vdd(vdd), .A(_3349_), .Y(_3350_) );
OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_3350_), .Y(_3351_) );
AOI21X1 AOI21X1_282 ( .gnd(gnd), .vdd(vdd), .A(_3348_), .B(_3350_), .C(_2005__bF_buf10), .Y(_3352_) );
AOI22X1 AOI22X1_801 ( .gnd(gnd), .vdd(vdd), .A(_2005__bF_buf9), .B(_3346_), .C(_3352_), .D(_3351_), .Y(_4__31_) );
NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf2), .B(_3375_), .Y(_3353_) );
OAI21X1 OAI21X1_1559 ( .gnd(gnd), .vdd(vdd), .A(_3375_), .B(_3387__bF_buf2), .C(_3353_), .Y(_11__0_) );
AOI22X1 AOI22X1_802 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf1), .B(_3377_), .C(round_ctr_reg_1_), .D(_113__bF_buf2), .Y(_3354_) );
AOI21X1 AOI21X1_283 ( .gnd(gnd), .vdd(vdd), .A(_3374_), .B(_3375_), .C(_3354_), .Y(_11__1_) );
INVX1 INVX1_1036 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_2_), .Y(_3355_) );
NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_2_), .B(_3376_), .Y(_3356_) );
AOI22X1 AOI22X1_803 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf0), .B(_3356_), .C(round_ctr_reg_2_), .D(_113__bF_buf1), .Y(_3357_) );
AOI21X1 AOI21X1_284 ( .gnd(gnd), .vdd(vdd), .A(_3355_), .B(_3377_), .C(_3357_), .Y(_11__2_) );
NOR2X1 NOR2X1_705 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_3380_), .Y(_3358_) );
INVX1 INVX1_1037 ( .gnd(gnd), .vdd(vdd), .A(_3358_), .Y(_3359_) );
OAI21X1 OAI21X1_1560 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf11), .B(_3370_), .C(round_ctr_reg_3_), .Y(_3360_) );
OAI21X1 OAI21X1_1561 ( .gnd(gnd), .vdd(vdd), .A(_3385_), .B(_3356_), .C(_3360_), .Y(_3361_) );
AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(_3359_), .B(_3361_), .Y(_11__3_) );
OAI21X1 OAI21X1_1562 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf10), .B(_3370_), .C(round_ctr_reg_4_), .Y(_3362_) );
MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_4_), .B(_3362_), .S(_3358_), .Y(_11__4_) );
INVX1 INVX1_1038 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_reg_4_), .Y(_3363_) );
OAI21X1 OAI21X1_1563 ( .gnd(gnd), .vdd(vdd), .A(_3363_), .B(_3380_), .C(_3400_), .Y(_3364_) );
OAI21X1 OAI21X1_1564 ( .gnd(gnd), .vdd(vdd), .A(_3380_), .B(_3389_), .C(_3364_), .Y(_3365_) );
OAI22X1 OAI22X1_133 ( .gnd(gnd), .vdd(vdd), .A(_3400_), .B(_3387__bF_buf1), .C(_3385_), .D(_3365_), .Y(_11__5_) );
NOR2X1 NOR2X1_706 ( .gnd(gnd), .vdd(vdd), .A(_3389_), .B(_3359_), .Y(_3366_) );
OAI21X1 OAI21X1_1565 ( .gnd(gnd), .vdd(vdd), .A(round_ctr_inc_bF_buf9), .B(_3370_), .C(round_ctr_reg_6_), .Y(_3367_) );
NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(_3388_), .B(_3366_), .Y(_3368_) );
OAI21X1 OAI21X1_1566 ( .gnd(gnd), .vdd(vdd), .A(_3366_), .B(_3367_), .C(_3368_), .Y(_11__6_) );
INVX1 INVX1_1039 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .Y(_3369_) );
OAI21X1 OAI21X1_1567 ( .gnd(gnd), .vdd(vdd), .A(_3369_), .B(round_ctr_rst_bF_buf60), .C(_2005__bF_buf8), .Y(_9_) );
NOR2X1 NOR2X1_707 ( .gnd(gnd), .vdd(vdd), .A(_3373_), .B(_3359_), .Y(_3665_) );
BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_3667__0_), .Y(digest[0]) );
BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_3667__1_), .Y(digest[1]) );
BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_3667__2_), .Y(digest[2]) );
BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_3667__3_), .Y(digest[3]) );
BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_3667__4_), .Y(digest[4]) );
BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_3667__5_), .Y(digest[5]) );
BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_3667__6_), .Y(digest[6]) );
BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_3667__7_), .Y(digest[7]) );
BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_3667__8_), .Y(digest[8]) );
BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_3667__9_), .Y(digest[9]) );
BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_3667__10_), .Y(digest[10]) );
BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_3667__11_), .Y(digest[11]) );
BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_3667__12_), .Y(digest[12]) );
BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_3667__13_), .Y(digest[13]) );
BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_3667__14_), .Y(digest[14]) );
BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_3667__15_), .Y(digest[15]) );
BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_3667__16_), .Y(digest[16]) );
BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_3667__17_), .Y(digest[17]) );
BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_3667__18_), .Y(digest[18]) );
BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_3667__19_), .Y(digest[19]) );
BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_3667__20_), .Y(digest[20]) );
BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_3667__21_), .Y(digest[21]) );
BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_3667__22_), .Y(digest[22]) );
BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_3667__23_), .Y(digest[23]) );
BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_3667__24_), .Y(digest[24]) );
BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_3667__25_), .Y(digest[25]) );
BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_3667__26_), .Y(digest[26]) );
BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_3667__27_), .Y(digest[27]) );
BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_3667__28_), .Y(digest[28]) );
BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_3667__29_), .Y(digest[29]) );
BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_3667__30_), .Y(digest[30]) );
BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(_3667__31_), .Y(digest[31]) );
BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(_3667__32_), .Y(digest[32]) );
BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(_3667__33_), .Y(digest[33]) );
BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(_3667__34_), .Y(digest[34]) );
BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(_3667__35_), .Y(digest[35]) );
BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(_3667__36_), .Y(digest[36]) );
BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(_3667__37_), .Y(digest[37]) );
BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(_3667__38_), .Y(digest[38]) );
BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(_3667__39_), .Y(digest[39]) );
BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(_3667__40_), .Y(digest[40]) );
BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(_3667__41_), .Y(digest[41]) );
BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(_3667__42_), .Y(digest[42]) );
BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(_3667__43_), .Y(digest[43]) );
BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(_3667__44_), .Y(digest[44]) );
BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(_3667__45_), .Y(digest[45]) );
BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(_3667__46_), .Y(digest[46]) );
BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(_3667__47_), .Y(digest[47]) );
BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(_3667__48_), .Y(digest[48]) );
BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(_3667__49_), .Y(digest[49]) );
BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(_3667__50_), .Y(digest[50]) );
BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(_3667__51_), .Y(digest[51]) );
BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(_3667__52_), .Y(digest[52]) );
BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(_3667__53_), .Y(digest[53]) );
BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(_3667__54_), .Y(digest[54]) );
BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(_3667__55_), .Y(digest[55]) );
BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(_3667__56_), .Y(digest[56]) );
BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(_3667__57_), .Y(digest[57]) );
BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(_3667__58_), .Y(digest[58]) );
BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(_3667__59_), .Y(digest[59]) );
BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(_3667__60_), .Y(digest[60]) );
BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(_3667__61_), .Y(digest[61]) );
BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(_3667__62_), .Y(digest[62]) );
BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(_3667__63_), .Y(digest[63]) );
BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(_3667__64_), .Y(digest[64]) );
BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(_3667__65_), .Y(digest[65]) );
BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(_3667__66_), .Y(digest[66]) );
BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(_3667__67_), .Y(digest[67]) );
BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(_3667__68_), .Y(digest[68]) );
BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(_3667__69_), .Y(digest[69]) );
BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(_3667__70_), .Y(digest[70]) );
BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(_3667__71_), .Y(digest[71]) );
BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(_3667__72_), .Y(digest[72]) );
BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(_3667__73_), .Y(digest[73]) );
BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(_3667__74_), .Y(digest[74]) );
BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(_3667__75_), .Y(digest[75]) );
BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(_3667__76_), .Y(digest[76]) );
BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(_3667__77_), .Y(digest[77]) );
BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(_3667__78_), .Y(digest[78]) );
BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(_3667__79_), .Y(digest[79]) );
BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(_3667__80_), .Y(digest[80]) );
BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(_3667__81_), .Y(digest[81]) );
BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(_3667__82_), .Y(digest[82]) );
BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(_3667__83_), .Y(digest[83]) );
BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(_3667__84_), .Y(digest[84]) );
BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(_3667__85_), .Y(digest[85]) );
BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(_3667__86_), .Y(digest[86]) );
BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(_3667__87_), .Y(digest[87]) );
BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(_3667__88_), .Y(digest[88]) );
BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(_3667__89_), .Y(digest[89]) );
BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(_3667__90_), .Y(digest[90]) );
BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(_3667__91_), .Y(digest[91]) );
BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(_3667__92_), .Y(digest[92]) );
BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(_3667__93_), .Y(digest[93]) );
BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(_3667__94_), .Y(digest[94]) );
BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(_3667__95_), .Y(digest[95]) );
BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(_3667__96_), .Y(digest[96]) );
BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(_3667__97_), .Y(digest[97]) );
BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(_3667__98_), .Y(digest[98]) );
BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(_3667__99_), .Y(digest[99]) );
BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(_3667__100_), .Y(digest[100]) );
BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(_3667__101_), .Y(digest[101]) );
BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(_3667__102_), .Y(digest[102]) );
BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(_3667__103_), .Y(digest[103]) );
BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(_3667__104_), .Y(digest[104]) );
BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(_3667__105_), .Y(digest[105]) );
BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(_3667__106_), .Y(digest[106]) );
BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(_3667__107_), .Y(digest[107]) );
BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(_3667__108_), .Y(digest[108]) );
BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(_3667__109_), .Y(digest[109]) );
BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(_3667__110_), .Y(digest[110]) );
BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(_3667__111_), .Y(digest[111]) );
BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(_3667__112_), .Y(digest[112]) );
BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(_3667__113_), .Y(digest[113]) );
BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(_3667__114_), .Y(digest[114]) );
BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(_3667__115_), .Y(digest[115]) );
BUFX2 BUFX2_127 ( .gnd(gnd), .vdd(vdd), .A(_3667__116_), .Y(digest[116]) );
BUFX2 BUFX2_128 ( .gnd(gnd), .vdd(vdd), .A(_3667__117_), .Y(digest[117]) );
BUFX2 BUFX2_129 ( .gnd(gnd), .vdd(vdd), .A(_3667__118_), .Y(digest[118]) );
BUFX2 BUFX2_130 ( .gnd(gnd), .vdd(vdd), .A(_3667__119_), .Y(digest[119]) );
BUFX2 BUFX2_131 ( .gnd(gnd), .vdd(vdd), .A(_3667__120_), .Y(digest[120]) );
BUFX2 BUFX2_132 ( .gnd(gnd), .vdd(vdd), .A(_3667__121_), .Y(digest[121]) );
BUFX2 BUFX2_133 ( .gnd(gnd), .vdd(vdd), .A(_3667__122_), .Y(digest[122]) );
BUFX2 BUFX2_134 ( .gnd(gnd), .vdd(vdd), .A(_3667__123_), .Y(digest[123]) );
BUFX2 BUFX2_135 ( .gnd(gnd), .vdd(vdd), .A(_3667__124_), .Y(digest[124]) );
BUFX2 BUFX2_136 ( .gnd(gnd), .vdd(vdd), .A(_3667__125_), .Y(digest[125]) );
BUFX2 BUFX2_137 ( .gnd(gnd), .vdd(vdd), .A(_3667__126_), .Y(digest[126]) );
BUFX2 BUFX2_138 ( .gnd(gnd), .vdd(vdd), .A(_3667__127_), .Y(digest[127]) );
BUFX2 BUFX2_139 ( .gnd(gnd), .vdd(vdd), .A(_3667__128_), .Y(digest[128]) );
BUFX2 BUFX2_140 ( .gnd(gnd), .vdd(vdd), .A(_3667__129_), .Y(digest[129]) );
BUFX2 BUFX2_141 ( .gnd(gnd), .vdd(vdd), .A(_3667__130_), .Y(digest[130]) );
BUFX2 BUFX2_142 ( .gnd(gnd), .vdd(vdd), .A(_3667__131_), .Y(digest[131]) );
BUFX2 BUFX2_143 ( .gnd(gnd), .vdd(vdd), .A(_3667__132_), .Y(digest[132]) );
BUFX2 BUFX2_144 ( .gnd(gnd), .vdd(vdd), .A(_3667__133_), .Y(digest[133]) );
BUFX2 BUFX2_145 ( .gnd(gnd), .vdd(vdd), .A(_3667__134_), .Y(digest[134]) );
BUFX2 BUFX2_146 ( .gnd(gnd), .vdd(vdd), .A(_3667__135_), .Y(digest[135]) );
BUFX2 BUFX2_147 ( .gnd(gnd), .vdd(vdd), .A(_3667__136_), .Y(digest[136]) );
BUFX2 BUFX2_148 ( .gnd(gnd), .vdd(vdd), .A(_3667__137_), .Y(digest[137]) );
BUFX2 BUFX2_149 ( .gnd(gnd), .vdd(vdd), .A(_3667__138_), .Y(digest[138]) );
BUFX2 BUFX2_150 ( .gnd(gnd), .vdd(vdd), .A(_3667__139_), .Y(digest[139]) );
BUFX2 BUFX2_151 ( .gnd(gnd), .vdd(vdd), .A(_3667__140_), .Y(digest[140]) );
BUFX2 BUFX2_152 ( .gnd(gnd), .vdd(vdd), .A(_3667__141_), .Y(digest[141]) );
BUFX2 BUFX2_153 ( .gnd(gnd), .vdd(vdd), .A(_3667__142_), .Y(digest[142]) );
BUFX2 BUFX2_154 ( .gnd(gnd), .vdd(vdd), .A(_3667__143_), .Y(digest[143]) );
BUFX2 BUFX2_155 ( .gnd(gnd), .vdd(vdd), .A(_3667__144_), .Y(digest[144]) );
BUFX2 BUFX2_156 ( .gnd(gnd), .vdd(vdd), .A(_3667__145_), .Y(digest[145]) );
BUFX2 BUFX2_157 ( .gnd(gnd), .vdd(vdd), .A(_3667__146_), .Y(digest[146]) );
BUFX2 BUFX2_158 ( .gnd(gnd), .vdd(vdd), .A(_3667__147_), .Y(digest[147]) );
BUFX2 BUFX2_159 ( .gnd(gnd), .vdd(vdd), .A(_3667__148_), .Y(digest[148]) );
BUFX2 BUFX2_160 ( .gnd(gnd), .vdd(vdd), .A(_3667__149_), .Y(digest[149]) );
BUFX2 BUFX2_161 ( .gnd(gnd), .vdd(vdd), .A(_3667__150_), .Y(digest[150]) );
BUFX2 BUFX2_162 ( .gnd(gnd), .vdd(vdd), .A(_3667__151_), .Y(digest[151]) );
BUFX2 BUFX2_163 ( .gnd(gnd), .vdd(vdd), .A(_3667__152_), .Y(digest[152]) );
BUFX2 BUFX2_164 ( .gnd(gnd), .vdd(vdd), .A(_3667__153_), .Y(digest[153]) );
BUFX2 BUFX2_165 ( .gnd(gnd), .vdd(vdd), .A(_3667__154_), .Y(digest[154]) );
BUFX2 BUFX2_166 ( .gnd(gnd), .vdd(vdd), .A(_3667__155_), .Y(digest[155]) );
BUFX2 BUFX2_167 ( .gnd(gnd), .vdd(vdd), .A(_3667__156_), .Y(digest[156]) );
BUFX2 BUFX2_168 ( .gnd(gnd), .vdd(vdd), .A(_3667__157_), .Y(digest[157]) );
BUFX2 BUFX2_169 ( .gnd(gnd), .vdd(vdd), .A(_3667__158_), .Y(digest[158]) );
BUFX2 BUFX2_170 ( .gnd(gnd), .vdd(vdd), .A(_3667__159_), .Y(digest[159]) );
BUFX2 BUFX2_171 ( .gnd(gnd), .vdd(vdd), .A(_3668_), .Y(digest_valid) );
BUFX2 BUFX2_172 ( .gnd(gnd), .vdd(vdd), .A(_3669_), .Y(ready) );
DFFSR DFFSR_514 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_3666__0_), .Q(_3669_), .R(vdd), .S(reset_n_bF_buf20) );
DFFSR DFFSR_515 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_3665_), .Q(digest_valid_new), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_516 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3666__2_), .Q(round_ctr_inc), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_517 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_5__0_), .Q(a_reg_0_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_518 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_5__1_), .Q(a_reg_1_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_519 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_5__2_), .Q(a_reg_2_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_520 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_5__3_), .Q(a_reg_3_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_521 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_5__4_), .Q(a_reg_4_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_522 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_5__5_), .Q(a_reg_5_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_523 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_5__6_), .Q(a_reg_6_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_524 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_5__7_), .Q(a_reg_7_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_525 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_5__8_), .Q(a_reg_8_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_526 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_5__9_), .Q(a_reg_9_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_527 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_5__10_), .Q(a_reg_10_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_528 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_5__11_), .Q(a_reg_11_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_529 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_5__12_), .Q(a_reg_12_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_530 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_5__13_), .Q(a_reg_13_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_531 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_5__14_), .Q(a_reg_14_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_532 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_5__15_), .Q(a_reg_15_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_533 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_5__16_), .Q(a_reg_16_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_534 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_5__17_), .Q(a_reg_17_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_535 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_5__18_), .Q(a_reg_18_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_536 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_5__19_), .Q(a_reg_19_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_537 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_5__20_), .Q(a_reg_20_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_538 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_5__21_), .Q(a_reg_21_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_539 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_5__22_), .Q(a_reg_22_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_540 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_5__23_), .Q(a_reg_23_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_541 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_5__24_), .Q(a_reg_24_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_542 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_5__25_), .Q(a_reg_25_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_543 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_5__26_), .Q(a_reg_26_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_544 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_5__27_), .Q(a_reg_27_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_545 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_5__28_), .Q(a_reg_28_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_546 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_5__29_), .Q(a_reg_29_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_547 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_5__30_), .Q(a_reg_30_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_548 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_5__31_), .Q(a_reg_31_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_549 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_6__0_), .Q(b_reg_0_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_550 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_6__1_), .Q(b_reg_1_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_551 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_6__2_), .Q(b_reg_2_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_552 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_6__3_), .Q(b_reg_3_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_553 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_6__4_), .Q(b_reg_4_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_554 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_6__5_), .Q(b_reg_5_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_555 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_6__6_), .Q(b_reg_6_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_556 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_6__7_), .Q(b_reg_7_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_557 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_6__8_), .Q(b_reg_8_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_558 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_6__9_), .Q(b_reg_9_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_559 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_6__10_), .Q(b_reg_10_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_560 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_6__11_), .Q(b_reg_11_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_561 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_6__12_), .Q(b_reg_12_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_562 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_6__13_), .Q(b_reg_13_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_563 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_6__14_), .Q(b_reg_14_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_564 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_6__15_), .Q(b_reg_15_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_565 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_6__16_), .Q(b_reg_16_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_566 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_6__17_), .Q(b_reg_17_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_567 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_6__18_), .Q(b_reg_18_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_568 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_6__19_), .Q(b_reg_19_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_569 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_6__20_), .Q(b_reg_20_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_570 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_6__21_), .Q(b_reg_21_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_571 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_6__22_), .Q(b_reg_22_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_572 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_6__23_), .Q(b_reg_23_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_573 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_6__24_), .Q(b_reg_24_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_574 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_6__25_), .Q(b_reg_25_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_575 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_6__26_), .Q(b_reg_26_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_576 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_6__27_), .Q(b_reg_27_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_577 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_6__28_), .Q(b_reg_28_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_578 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_6__29_), .Q(b_reg_29_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_579 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_6__30_), .Q(b_reg_30_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_580 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_6__31_), .Q(b_reg_31_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_581 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_7__0_), .Q(c_reg_0_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_582 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_7__1_), .Q(c_reg_1_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_583 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_7__2_), .Q(c_reg_2_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_584 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_7__3_), .Q(c_reg_3_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_585 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_7__4_), .Q(c_reg_4_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_586 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_7__5_), .Q(c_reg_5_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_587 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_7__6_), .Q(c_reg_6_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_588 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_7__7_), .Q(c_reg_7_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_589 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_7__8_), .Q(c_reg_8_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_590 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_7__9_), .Q(c_reg_9_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_591 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_7__10_), .Q(c_reg_10_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_592 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_7__11_), .Q(c_reg_11_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_593 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_7__12_), .Q(c_reg_12_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_594 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_7__13_), .Q(c_reg_13_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_595 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_7__14_), .Q(c_reg_14_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_596 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_7__15_), .Q(c_reg_15_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_597 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_7__16_), .Q(c_reg_16_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_598 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_7__17_), .Q(c_reg_17_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_599 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_7__18_), .Q(c_reg_18_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_600 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_7__19_), .Q(c_reg_19_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_601 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_7__20_), .Q(c_reg_20_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_602 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_7__21_), .Q(c_reg_21_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_603 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_7__22_), .Q(c_reg_22_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_604 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_7__23_), .Q(c_reg_23_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_605 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_7__24_), .Q(c_reg_24_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_606 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_7__25_), .Q(c_reg_25_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_607 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_7__26_), .Q(c_reg_26_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_608 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_7__27_), .Q(c_reg_27_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_609 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_7__28_), .Q(c_reg_28_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_610 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_7__29_), .Q(c_reg_29_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_611 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_7__30_), .Q(c_reg_30_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_612 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_7__31_), .Q(c_reg_31_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_613 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_8__0_), .Q(d_reg_0_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_614 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_8__1_), .Q(d_reg_1_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_615 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_8__2_), .Q(d_reg_2_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_616 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_8__3_), .Q(d_reg_3_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_617 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_8__4_), .Q(d_reg_4_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_618 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_8__5_), .Q(d_reg_5_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_619 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_8__6_), .Q(d_reg_6_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_620 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_8__7_), .Q(d_reg_7_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_621 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_8__8_), .Q(d_reg_8_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_622 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_8__9_), .Q(d_reg_9_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_623 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_8__10_), .Q(d_reg_10_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_624 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_8__11_), .Q(d_reg_11_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_625 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_8__12_), .Q(d_reg_12_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_626 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_8__13_), .Q(d_reg_13_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_627 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_8__14_), .Q(d_reg_14_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_628 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_8__15_), .Q(d_reg_15_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_629 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_8__16_), .Q(d_reg_16_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_630 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_8__17_), .Q(d_reg_17_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_631 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_8__18_), .Q(d_reg_18_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_632 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_8__19_), .Q(d_reg_19_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_633 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_8__20_), .Q(d_reg_20_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_634 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_8__21_), .Q(d_reg_21_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_635 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_8__22_), .Q(d_reg_22_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_636 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_8__23_), .Q(d_reg_23_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_637 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_8__24_), .Q(d_reg_24_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_638 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_8__25_), .Q(d_reg_25_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_639 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_8__26_), .Q(d_reg_26_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_640 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_8__27_), .Q(d_reg_27_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_641 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_8__28_), .Q(d_reg_28_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_642 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_8__29_), .Q(d_reg_29_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_643 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_8__30_), .Q(d_reg_30_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_644 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_8__31_), .Q(d_reg_31_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_645 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_10__0_), .Q(e_reg_0_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_646 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_10__1_), .Q(e_reg_1_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_647 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_10__2_), .Q(e_reg_2_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_648 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_10__3_), .Q(e_reg_3_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_649 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_10__4_), .Q(e_reg_4_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_650 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_10__5_), .Q(e_reg_5_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_651 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_10__6_), .Q(e_reg_6_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_652 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_10__7_), .Q(e_reg_7_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_653 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_10__8_), .Q(e_reg_8_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_654 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_10__9_), .Q(e_reg_9_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_655 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_10__10_), .Q(e_reg_10_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_656 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_10__11_), .Q(e_reg_11_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_657 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_10__12_), .Q(e_reg_12_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_658 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_10__13_), .Q(e_reg_13_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_659 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_10__14_), .Q(e_reg_14_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_660 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_10__15_), .Q(e_reg_15_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_661 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_10__16_), .Q(e_reg_16_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_662 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_10__17_), .Q(e_reg_17_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_663 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_10__18_), .Q(e_reg_18_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_664 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_10__19_), .Q(e_reg_19_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_665 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_10__20_), .Q(e_reg_20_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_666 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_10__21_), .Q(e_reg_21_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_667 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_10__22_), .Q(e_reg_22_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_668 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_10__23_), .Q(e_reg_23_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_669 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_10__24_), .Q(e_reg_24_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_670 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_10__25_), .Q(e_reg_25_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_671 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_10__26_), .Q(e_reg_26_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_672 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_10__27_), .Q(e_reg_27_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_673 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_10__28_), .Q(e_reg_28_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_674 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_10__29_), .Q(e_reg_29_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_675 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_10__30_), .Q(e_reg_30_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_676 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_10__31_), .Q(e_reg_31_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_677 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_0__0_), .Q(_3667__128_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_678 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_0__1_), .Q(_3667__129_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_679 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_0__2_), .Q(_3667__130_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_680 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_0__3_), .Q(_3667__131_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_681 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_0__4_), .Q(_3667__132_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_682 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_0__5_), .Q(_3667__133_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_683 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_0__6_), .Q(_3667__134_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_684 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_0__7_), .Q(_3667__135_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_685 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_0__8_), .Q(_3667__136_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_686 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_0__9_), .Q(_3667__137_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_687 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_0__10_), .Q(_3667__138_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_688 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_0__11_), .Q(_3667__139_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_689 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_0__12_), .Q(_3667__140_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_690 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_0__13_), .Q(_3667__141_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_691 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_0__14_), .Q(_3667__142_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_692 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_0__15_), .Q(_3667__143_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_693 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_0__16_), .Q(_3667__144_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_694 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_0__17_), .Q(_3667__145_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_695 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_0__18_), .Q(_3667__146_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_696 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_0__19_), .Q(_3667__147_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_697 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_0__20_), .Q(_3667__148_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_698 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_0__21_), .Q(_3667__149_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_699 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0__22_), .Q(_3667__150_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_700 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__23_), .Q(_3667__151_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_701 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__24_), .Q(_3667__152_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_702 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__25_), .Q(_3667__153_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_703 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__26_), .Q(_3667__154_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_704 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__27_), .Q(_3667__155_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_705 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__28_), .Q(_3667__156_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_706 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_0__29_), .Q(_3667__157_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_707 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_0__30_), .Q(_3667__158_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_708 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_0__31_), .Q(_3667__159_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_709 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_1__0_), .Q(_3667__96_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_710 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_1__1_), .Q(_3667__97_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_711 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_1__2_), .Q(_3667__98_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_712 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_1__3_), .Q(_3667__99_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_713 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_1__4_), .Q(_3667__100_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_714 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_1__5_), .Q(_3667__101_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_715 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_1__6_), .Q(_3667__102_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_716 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_1__7_), .Q(_3667__103_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_717 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_1__8_), .Q(_3667__104_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_718 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_1__9_), .Q(_3667__105_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_719 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_1__10_), .Q(_3667__106_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_720 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_1__11_), .Q(_3667__107_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_721 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_1__12_), .Q(_3667__108_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_722 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_1__13_), .Q(_3667__109_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_723 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_1__14_), .Q(_3667__110_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_724 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_1__15_), .Q(_3667__111_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_725 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_1__16_), .Q(_3667__112_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_726 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_1__17_), .Q(_3667__113_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_727 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_1__18_), .Q(_3667__114_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_728 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_1__19_), .Q(_3667__115_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_729 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_1__20_), .Q(_3667__116_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_730 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_1__21_), .Q(_3667__117_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_731 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_1__22_), .Q(_3667__118_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_732 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_1__23_), .Q(_3667__119_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_733 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_1__24_), .Q(_3667__120_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_734 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_1__25_), .Q(_3667__121_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_735 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_1__26_), .Q(_3667__122_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_736 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_1__27_), .Q(_3667__123_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_737 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_1__28_), .Q(_3667__124_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_738 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_1768_), .Q(_3667__125_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_739 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_1__30_), .Q(_3667__126_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_740 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_1__31_), .Q(_3667__127_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_741 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_2__0_), .Q(_3667__64_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_742 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_2__1_), .Q(_3667__65_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_743 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_2__2_), .Q(_3667__66_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_744 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_2__3_), .Q(_3667__67_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_745 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_2__4_), .Q(_3667__68_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_746 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_2__5_), .Q(_3667__69_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_747 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_2__6_), .Q(_3667__70_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_748 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_2__7_), .Q(_3667__71_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_749 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_2__8_), .Q(_3667__72_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_750 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_2__9_), .Q(_3667__73_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_751 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_2__10_), .Q(_3667__74_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_752 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_2__11_), .Q(_3667__75_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_753 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_2__12_), .Q(_3667__76_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_754 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_2__13_), .Q(_3667__77_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_755 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_2__14_), .Q(_3667__78_), .R(reset_n_bF_buf46), .S(vdd) );
DFFSR DFFSR_756 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf38), .D(_2__15_), .Q(_3667__79_), .R(reset_n_bF_buf45), .S(vdd) );
DFFSR DFFSR_757 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf37), .D(_2__16_), .Q(_3667__80_), .R(reset_n_bF_buf44), .S(vdd) );
DFFSR DFFSR_758 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf36), .D(_2__17_), .Q(_3667__81_), .R(reset_n_bF_buf43), .S(vdd) );
DFFSR DFFSR_759 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf35), .D(_2__18_), .Q(_3667__82_), .R(reset_n_bF_buf42), .S(vdd) );
DFFSR DFFSR_760 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf34), .D(_2__19_), .Q(_3667__83_), .R(reset_n_bF_buf41), .S(vdd) );
DFFSR DFFSR_761 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf33), .D(_2__20_), .Q(_3667__84_), .R(reset_n_bF_buf40), .S(vdd) );
DFFSR DFFSR_762 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf32), .D(_2__21_), .Q(_3667__85_), .R(reset_n_bF_buf39), .S(vdd) );
DFFSR DFFSR_763 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf31), .D(_2__22_), .Q(_3667__86_), .R(reset_n_bF_buf38), .S(vdd) );
DFFSR DFFSR_764 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf30), .D(_2__23_), .Q(_3667__87_), .R(reset_n_bF_buf37), .S(vdd) );
DFFSR DFFSR_765 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf29), .D(_2__24_), .Q(_3667__88_), .R(reset_n_bF_buf36), .S(vdd) );
DFFSR DFFSR_766 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf28), .D(_2__25_), .Q(_3667__89_), .R(reset_n_bF_buf35), .S(vdd) );
DFFSR DFFSR_767 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf27), .D(_2__26_), .Q(_3667__90_), .R(reset_n_bF_buf34), .S(vdd) );
DFFSR DFFSR_768 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf26), .D(_2__27_), .Q(_3667__91_), .R(reset_n_bF_buf33), .S(vdd) );
DFFSR DFFSR_769 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf25), .D(_2__28_), .Q(_3667__92_), .R(reset_n_bF_buf32), .S(vdd) );
DFFSR DFFSR_770 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf24), .D(_2__29_), .Q(_3667__93_), .R(reset_n_bF_buf31), .S(vdd) );
DFFSR DFFSR_771 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf23), .D(_2__30_), .Q(_3667__94_), .R(reset_n_bF_buf30), .S(vdd) );
DFFSR DFFSR_772 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf22), .D(_2__31_), .Q(_3667__95_), .R(reset_n_bF_buf29), .S(vdd) );
DFFSR DFFSR_773 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf21), .D(_3__0_), .Q(_3667__32_), .R(reset_n_bF_buf28), .S(vdd) );
DFFSR DFFSR_774 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf20), .D(_3__1_), .Q(_3667__33_), .R(reset_n_bF_buf27), .S(vdd) );
DFFSR DFFSR_775 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf19), .D(_3__2_), .Q(_3667__34_), .R(reset_n_bF_buf26), .S(vdd) );
DFFSR DFFSR_776 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf18), .D(_3__3_), .Q(_3667__35_), .R(reset_n_bF_buf25), .S(vdd) );
DFFSR DFFSR_777 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf17), .D(_3__4_), .Q(_3667__36_), .R(reset_n_bF_buf24), .S(vdd) );
DFFSR DFFSR_778 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf16), .D(_3__5_), .Q(_3667__37_), .R(reset_n_bF_buf23), .S(vdd) );
DFFSR DFFSR_779 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf15), .D(_3__6_), .Q(_3667__38_), .R(reset_n_bF_buf22), .S(vdd) );
DFFSR DFFSR_780 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf14), .D(_3__7_), .Q(_3667__39_), .R(reset_n_bF_buf21), .S(vdd) );
DFFSR DFFSR_781 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf13), .D(_3__8_), .Q(_3667__40_), .R(reset_n_bF_buf20), .S(vdd) );
DFFSR DFFSR_782 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf12), .D(_3__9_), .Q(_3667__41_), .R(reset_n_bF_buf19), .S(vdd) );
DFFSR DFFSR_783 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf11), .D(_3__10_), .Q(_3667__42_), .R(reset_n_bF_buf18), .S(vdd) );
DFFSR DFFSR_784 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf10), .D(_3__11_), .Q(_3667__43_), .R(reset_n_bF_buf17), .S(vdd) );
DFFSR DFFSR_785 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf9), .D(_3__12_), .Q(_3667__44_), .R(reset_n_bF_buf16), .S(vdd) );
DFFSR DFFSR_786 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_3__13_), .Q(_3667__45_), .R(reset_n_bF_buf15), .S(vdd) );
DFFSR DFFSR_787 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_3__14_), .Q(_3667__46_), .R(reset_n_bF_buf14), .S(vdd) );
DFFSR DFFSR_788 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_3__15_), .Q(_3667__47_), .R(reset_n_bF_buf13), .S(vdd) );
DFFSR DFFSR_789 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_3__16_), .Q(_3667__48_), .R(reset_n_bF_buf12), .S(vdd) );
DFFSR DFFSR_790 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3__17_), .Q(_3667__49_), .R(reset_n_bF_buf11), .S(vdd) );
DFFSR DFFSR_791 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_3__18_), .Q(_3667__50_), .R(reset_n_bF_buf10), .S(vdd) );
DFFSR DFFSR_792 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_3__19_), .Q(_3667__51_), .R(reset_n_bF_buf9), .S(vdd) );
DFFSR DFFSR_793 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_3__20_), .Q(_3667__52_), .R(reset_n_bF_buf8), .S(vdd) );
DFFSR DFFSR_794 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_3__21_), .Q(_3667__53_), .R(reset_n_bF_buf7), .S(vdd) );
DFFSR DFFSR_795 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf88), .D(_3__22_), .Q(_3667__54_), .R(reset_n_bF_buf6), .S(vdd) );
DFFSR DFFSR_796 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf87), .D(_3__23_), .Q(_3667__55_), .R(reset_n_bF_buf5), .S(vdd) );
DFFSR DFFSR_797 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf86), .D(_3__24_), .Q(_3667__56_), .R(reset_n_bF_buf4), .S(vdd) );
DFFSR DFFSR_798 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf85), .D(_3__25_), .Q(_3667__57_), .R(reset_n_bF_buf3), .S(vdd) );
DFFSR DFFSR_799 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf84), .D(_3__26_), .Q(_3667__58_), .R(reset_n_bF_buf2), .S(vdd) );
DFFSR DFFSR_800 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf83), .D(_3__27_), .Q(_3667__59_), .R(reset_n_bF_buf1), .S(vdd) );
DFFSR DFFSR_801 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf82), .D(_3__28_), .Q(_3667__60_), .R(reset_n_bF_buf0), .S(vdd) );
DFFSR DFFSR_802 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf81), .D(_3__29_), .Q(_3667__61_), .R(reset_n_bF_buf88), .S(vdd) );
DFFSR DFFSR_803 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf80), .D(_3__30_), .Q(_3667__62_), .R(reset_n_bF_buf87), .S(vdd) );
DFFSR DFFSR_804 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf79), .D(_3__31_), .Q(_3667__63_), .R(reset_n_bF_buf86), .S(vdd) );
DFFSR DFFSR_805 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf78), .D(_4__0_), .Q(_3667__0_), .R(reset_n_bF_buf85), .S(vdd) );
DFFSR DFFSR_806 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf77), .D(_4__1_), .Q(_3667__1_), .R(reset_n_bF_buf84), .S(vdd) );
DFFSR DFFSR_807 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf76), .D(_4__2_), .Q(_3667__2_), .R(reset_n_bF_buf83), .S(vdd) );
DFFSR DFFSR_808 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf75), .D(_4__3_), .Q(_3667__3_), .R(reset_n_bF_buf82), .S(vdd) );
DFFSR DFFSR_809 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf74), .D(_4__4_), .Q(_3667__4_), .R(reset_n_bF_buf81), .S(vdd) );
DFFSR DFFSR_810 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf73), .D(_4__5_), .Q(_3667__5_), .R(reset_n_bF_buf80), .S(vdd) );
DFFSR DFFSR_811 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf72), .D(_4__6_), .Q(_3667__6_), .R(reset_n_bF_buf79), .S(vdd) );
DFFSR DFFSR_812 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf71), .D(_4__7_), .Q(_3667__7_), .R(reset_n_bF_buf78), .S(vdd) );
DFFSR DFFSR_813 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf70), .D(_4__8_), .Q(_3667__8_), .R(reset_n_bF_buf77), .S(vdd) );
DFFSR DFFSR_814 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf69), .D(_4__9_), .Q(_3667__9_), .R(reset_n_bF_buf76), .S(vdd) );
DFFSR DFFSR_815 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf68), .D(_4__10_), .Q(_3667__10_), .R(reset_n_bF_buf75), .S(vdd) );
DFFSR DFFSR_816 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf67), .D(_4__11_), .Q(_3667__11_), .R(reset_n_bF_buf74), .S(vdd) );
DFFSR DFFSR_817 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf66), .D(_4__12_), .Q(_3667__12_), .R(reset_n_bF_buf73), .S(vdd) );
DFFSR DFFSR_818 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf65), .D(_4__13_), .Q(_3667__13_), .R(reset_n_bF_buf72), .S(vdd) );
DFFSR DFFSR_819 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf64), .D(_4__14_), .Q(_3667__14_), .R(reset_n_bF_buf71), .S(vdd) );
DFFSR DFFSR_820 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf63), .D(_4__15_), .Q(_3667__15_), .R(reset_n_bF_buf70), .S(vdd) );
DFFSR DFFSR_821 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf62), .D(_4__16_), .Q(_3667__16_), .R(reset_n_bF_buf69), .S(vdd) );
DFFSR DFFSR_822 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf61), .D(_4__17_), .Q(_3667__17_), .R(reset_n_bF_buf68), .S(vdd) );
DFFSR DFFSR_823 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf60), .D(_4__18_), .Q(_3667__18_), .R(reset_n_bF_buf67), .S(vdd) );
DFFSR DFFSR_824 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf59), .D(_4__19_), .Q(_3667__19_), .R(reset_n_bF_buf66), .S(vdd) );
DFFSR DFFSR_825 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf58), .D(_4__20_), .Q(_3667__20_), .R(reset_n_bF_buf65), .S(vdd) );
DFFSR DFFSR_826 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf57), .D(_4__21_), .Q(_3667__21_), .R(reset_n_bF_buf64), .S(vdd) );
DFFSR DFFSR_827 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf56), .D(_4__22_), .Q(_3667__22_), .R(reset_n_bF_buf63), .S(vdd) );
DFFSR DFFSR_828 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf55), .D(_4__23_), .Q(_3667__23_), .R(reset_n_bF_buf62), .S(vdd) );
DFFSR DFFSR_829 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf54), .D(_4__24_), .Q(_3667__24_), .R(reset_n_bF_buf61), .S(vdd) );
DFFSR DFFSR_830 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf53), .D(_4__25_), .Q(_3667__25_), .R(reset_n_bF_buf60), .S(vdd) );
DFFSR DFFSR_831 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf52), .D(_4__26_), .Q(_3667__26_), .R(reset_n_bF_buf59), .S(vdd) );
DFFSR DFFSR_832 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf51), .D(_4__27_), .Q(_3667__27_), .R(reset_n_bF_buf58), .S(vdd) );
DFFSR DFFSR_833 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf50), .D(_4__28_), .Q(_3667__28_), .R(reset_n_bF_buf57), .S(vdd) );
DFFSR DFFSR_834 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf49), .D(_4__29_), .Q(_3667__29_), .R(reset_n_bF_buf56), .S(vdd) );
DFFSR DFFSR_835 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf48), .D(_4__30_), .Q(_3667__30_), .R(reset_n_bF_buf55), .S(vdd) );
DFFSR DFFSR_836 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf47), .D(_4__31_), .Q(_3667__31_), .R(reset_n_bF_buf54), .S(vdd) );
DFFSR DFFSR_837 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf46), .D(_11__0_), .Q(round_ctr_reg_0_), .R(reset_n_bF_buf53), .S(vdd) );
DFFSR DFFSR_838 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf45), .D(_11__1_), .Q(round_ctr_reg_1_), .R(reset_n_bF_buf52), .S(vdd) );
DFFSR DFFSR_839 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf44), .D(_11__2_), .Q(round_ctr_reg_2_), .R(reset_n_bF_buf51), .S(vdd) );
DFFSR DFFSR_840 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf43), .D(_11__3_), .Q(round_ctr_reg_3_), .R(reset_n_bF_buf50), .S(vdd) );
DFFSR DFFSR_841 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf42), .D(_11__4_), .Q(round_ctr_reg_4_), .R(reset_n_bF_buf49), .S(vdd) );
DFFSR DFFSR_842 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf41), .D(_11__5_), .Q(round_ctr_reg_5_), .R(reset_n_bF_buf48), .S(vdd) );
DFFSR DFFSR_843 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf40), .D(_11__6_), .Q(round_ctr_reg_6_), .R(reset_n_bF_buf47), .S(vdd) );
DFFSR DFFSR_844 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf39), .D(_9_), .Q(_3668_), .R(reset_n_bF_buf46), .S(vdd) );
INVX1 INVX1_1040 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_4_), .Y(_3688_) );
INVX1 INVX1_1041 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_5_), .Y(_3689_) );
NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(_3688_), .B(_3689_), .Y(_3690_) );
NOR2X1 NOR2X1_708 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_6_), .B(_3690_), .Y(_3691_) );
INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(_3691__bF_buf0), .Y(_3692_) );
XNOR2X1 XNOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__31_), .B(w_mem_inst_w_mem_8__31_), .Y(_3693_) );
XNOR2X1 XNOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst_w_mem_0__31_), .Y(_3694_) );
XNOR2X1 XNOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(_3693_), .B(_3694_), .Y(_3695_) );
INVX1 INVX1_1042 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__0_), .Y(_3696_) );
OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .Y(_3697_) );
INVX2 INVX2_85 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_0_), .Y(_3698_) );
NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_1_), .B(_3698_), .Y(_3699_) );
NOR2X1 NOR2X1_709 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3699_), .Y(_3700_) );
INVX4 INVX4_6 ( .gnd(gnd), .vdd(vdd), .A(_3700__bF_buf3), .Y(_3701_) );
OAI21X1 OAI21X1_1568 ( .gnd(gnd), .vdd(vdd), .A(_3696_), .B(_3701_), .C(_3691__bF_buf4), .Y(_3702_) );
INVX1 INVX1_1043 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__0_), .Y(_3703_) );
INVX1 INVX1_1044 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_3_), .Y(_3704_) );
NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_2_), .B(_3704_), .Y(_3705_) );
NOR2X1 NOR2X1_710 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3705_), .Y(_3706_) );
INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(_3706__bF_buf3), .Y(_3707_) );
NOR2X1 NOR2X1_711 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(_3708_) );
NOR2X1 NOR2X1_712 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .Y(_3709_) );
AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(_3708_), .B(_3709_), .Y(_3710_) );
NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__0_), .B(_3710__bF_buf0), .Y(_3711_) );
OAI21X1 OAI21X1_1569 ( .gnd(gnd), .vdd(vdd), .A(_3703_), .B(_3707_), .C(_3711_), .Y(_3712_) );
INVX1 INVX1_1045 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__0_), .Y(_3713_) );
INVX1 INVX1_1046 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__0_), .Y(_3714_) );
NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .Y(_3715_) );
NOR3X1 NOR3X1_86 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_1_), .B(_3698_), .C(_3715_), .Y(_3716_) );
INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .Y(_3717_) );
OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(_3718_) );
INVX2 INVX2_86 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_2_), .Y(_3719_) );
NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_3_), .B(_3719_), .Y(_3720_) );
NOR2X1 NOR2X1_713 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .B(_3720_), .Y(_3721_) );
INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(_3721_), .Y(_3722_) );
OAI22X1 OAI22X1_134 ( .gnd(gnd), .vdd(vdd), .A(_3714_), .B(_3717__bF_buf1), .C(_3713_), .D(_3722__bF_buf3), .Y(_3723_) );
NOR3X1 NOR3X1_87 ( .gnd(gnd), .vdd(vdd), .A(_3702_), .B(_3723_), .C(_3712_), .Y(_3724_) );
INVX2 INVX2_87 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_1_), .Y(_3725_) );
NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_0_), .B(_3725_), .Y(_3726_) );
NOR2X1 NOR2X1_714 ( .gnd(gnd), .vdd(vdd), .A(_3726_), .B(_3720_), .Y(_3727_) );
NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__0_), .B(_3727__bF_buf1), .Y(_3728_) );
NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(_3729_) );
NOR2X1 NOR2X1_715 ( .gnd(gnd), .vdd(vdd), .A(_3729_), .B(_3697_), .Y(_3730_) );
NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__0_), .B(_3730__bF_buf2), .Y(_3731_) );
NOR2X1 NOR2X1_716 ( .gnd(gnd), .vdd(vdd), .A(_3697_), .B(_3726_), .Y(_3732_) );
NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__0_), .B(_3732__bF_buf1), .Y(_3733_) );
NAND3X1 NAND3X1_312 ( .gnd(gnd), .vdd(vdd), .A(_3731_), .B(_3733_), .C(_3728_), .Y(_3734_) );
NOR3X1 NOR3X1_88 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_0_), .B(_3725_), .C(_3715_), .Y(_3735_) );
NOR3X1 NOR3X1_89 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_3_), .B(_3719_), .C(_3729_), .Y(_3736_) );
AOI22X1 AOI22X1_804 ( .gnd(gnd), .vdd(vdd), .A(_3735__bF_buf0), .B(w_mem_inst_w_mem_14__0_), .C(w_mem_inst_w_mem_7__0_), .D(_3736__bF_buf0), .Y(_3737_) );
NOR2X1 NOR2X1_717 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_3729_), .Y(_3738_) );
NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__0_), .B(_3738__bF_buf3), .Y(_3739_) );
NOR2X1 NOR2X1_718 ( .gnd(gnd), .vdd(vdd), .A(_3718_), .B(_3705_), .Y(_3740_) );
NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__0_), .B(_3740__bF_buf0), .Y(_3741_) );
NAND3X1 NAND3X1_313 ( .gnd(gnd), .vdd(vdd), .A(_3739_), .B(_3741_), .C(_3737_), .Y(_3742_) );
NOR2X1 NOR2X1_719 ( .gnd(gnd), .vdd(vdd), .A(_3705_), .B(_3726_), .Y(_3743_) );
NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__0_), .B(_3743_), .Y(_3744_) );
NOR3X1 NOR3X1_90 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_ctr_reg_2_), .B(_3704_), .C(_3729_), .Y(_3745_) );
NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__0_), .B(_3745__bF_buf0), .Y(_3746_) );
NOR2X1 NOR2X1_720 ( .gnd(gnd), .vdd(vdd), .A(_3715_), .B(_3718_), .Y(_3747_) );
NOR2X1 NOR2X1_721 ( .gnd(gnd), .vdd(vdd), .A(_3699_), .B(_3720_), .Y(_3748_) );
AOI22X1 AOI22X1_805 ( .gnd(gnd), .vdd(vdd), .A(_3747__bF_buf0), .B(w_mem_inst_w_mem_12__0_), .C(w_mem_inst_w_mem_10__0_), .D(_3748__bF_buf4), .Y(_3749_) );
NAND3X1 NAND3X1_314 ( .gnd(gnd), .vdd(vdd), .A(_3744_), .B(_3746_), .C(_3749_), .Y(_3750_) );
NOR3X1 NOR3X1_91 ( .gnd(gnd), .vdd(vdd), .A(_3734_), .B(_3742_), .C(_3750_), .Y(_3751_) );
AOI22X1 AOI22X1_806 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf4), .B(_3695_), .C(_3724_), .D(_3751_), .Y(w_0_) );
XNOR2X1 XNOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__0_), .B(w_mem_inst_w_mem_13__0_), .Y(_3752_) );
XNOR2X1 XNOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__0_), .B(w_mem_inst_w_mem_2__0_), .Y(_3753_) );
XNOR2X1 XNOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(_3752_), .B(_3753_), .Y(_3754_) );
INVX1 INVX1_1047 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__1_), .Y(_3755_) );
OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(_3705_), .B(_3726_), .Y(_3756_) );
OAI21X1 OAI21X1_1570 ( .gnd(gnd), .vdd(vdd), .A(_3755_), .B(_3756_), .C(_3691__bF_buf3), .Y(_3757_) );
INVX1 INVX1_1048 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_13__1_), .Y(_3758_) );
NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__1_), .B(_3747__bF_buf4), .Y(_3759_) );
OAI21X1 OAI21X1_1571 ( .gnd(gnd), .vdd(vdd), .A(_3758_), .B(_3717__bF_buf0), .C(_3759_), .Y(_3760_) );
INVX1 INVX1_1049 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__1_), .Y(_3761_) );
INVX1 INVX1_1050 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__1_), .Y(_3762_) );
INVX4 INVX4_7 ( .gnd(gnd), .vdd(vdd), .A(_3727__bF_buf0), .Y(_3763_) );
INVX4 INVX4_8 ( .gnd(gnd), .vdd(vdd), .A(_3730__bF_buf1), .Y(_3764_) );
OAI22X1 OAI22X1_135 ( .gnd(gnd), .vdd(vdd), .A(_3762_), .B(_3764_), .C(_3761_), .D(_3763_), .Y(_3765_) );
NOR3X1 NOR3X1_92 ( .gnd(gnd), .vdd(vdd), .A(_3757_), .B(_3760_), .C(_3765_), .Y(_3766_) );
NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__1_), .B(_3738__bF_buf2), .Y(_3767_) );
NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_4__1_), .B(_3740__bF_buf3), .Y(_3768_) );
NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__1_), .B(_3710__bF_buf4), .Y(_3769_) );
NAND3X1 NAND3X1_315 ( .gnd(gnd), .vdd(vdd), .A(_3767_), .B(_3769_), .C(_3768_), .Y(_3770_) );
AOI22X1 AOI22X1_807 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_7__1_), .B(_3736__bF_buf3), .C(w_mem_inst_w_mem_2__1_), .D(_3700__bF_buf2), .Y(_3771_) );
AOI22X1 AOI22X1_808 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__1_), .B(_3745__bF_buf4), .C(w_mem_inst_w_mem_1__1_), .D(_3732__bF_buf0), .Y(_3772_) );
NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(_3771_), .B(_3772_), .Y(_3773_) );
AOI22X1 AOI22X1_809 ( .gnd(gnd), .vdd(vdd), .A(_3721_), .B(w_mem_inst_w_mem_8__1_), .C(w_mem_inst_w_mem_6__1_), .D(_3706__bF_buf2), .Y(_3774_) );
NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_14__1_), .B(_3735__bF_buf4), .Y(_3775_) );
NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__1_), .B(_3748__bF_buf3), .Y(_3776_) );
NAND3X1 NAND3X1_316 ( .gnd(gnd), .vdd(vdd), .A(_3775_), .B(_3776_), .C(_3774_), .Y(_3777_) );
NOR3X1 NOR3X1_93 ( .gnd(gnd), .vdd(vdd), .A(_3770_), .B(_3773_), .C(_3777_), .Y(_3778_) );
AOI22X1 AOI22X1_810 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf3), .B(_3754_), .C(_3766_), .D(_3778_), .Y(w_1_) );
XNOR2X1 XNOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__1_), .B(w_mem_inst_w_mem_13__1_), .Y(_3779_) );
XNOR2X1 XNOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__1_), .B(w_mem_inst_w_mem_2__1_), .Y(_3780_) );
XNOR2X1 XNOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(_3779_), .B(_3780_), .Y(_3781_) );
INVX1 INVX1_1051 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_10__2_), .Y(_3782_) );
INVX2 INVX2_88 ( .gnd(gnd), .vdd(vdd), .A(_3748__bF_buf2), .Y(_3783_) );
OAI21X1 OAI21X1_1572 ( .gnd(gnd), .vdd(vdd), .A(_3782_), .B(_3783_), .C(_3691__bF_buf2), .Y(_3784_) );
INVX1 INVX1_1052 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_9__2_), .Y(_3785_) );
NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_12__2_), .B(_3747__bF_buf3), .Y(_3786_) );
OAI21X1 OAI21X1_1573 ( .gnd(gnd), .vdd(vdd), .A(_3785_), .B(_3763_), .C(_3786_), .Y(_3787_) );
INVX1 INVX1_1053 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_1__2_), .Y(_3788_) );
INVX1 INVX1_1054 ( .gnd(gnd), .vdd(vdd), .A(_3732__bF_buf4), .Y(_3789_) );
NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__2_), .B(_3710__bF_buf3), .Y(_3790_) );
OAI21X1 OAI21X1_1574 ( .gnd(gnd), .vdd(vdd), .A(_3788_), .B(_3789_), .C(_3790_), .Y(_3791_) );
NOR3X1 NOR3X1_94 ( .gnd(gnd), .vdd(vdd), .A(_3791_), .B(_3784_), .C(_3787_), .Y(_3792_) );
INVX1 INVX1_1055 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_5__2_), .Y(_3793_) );
AOI22X1 AOI22X1_811 ( .gnd(gnd), .vdd(vdd), .A(_3716_), .B(w_mem_inst_w_mem_13__2_), .C(w_mem_inst_w_mem_14__2_), .D(_3735__bF_buf3), .Y(_3794_) );
OAI21X1 OAI21X1_1575 ( .gnd(gnd), .vdd(vdd), .A(_3793_), .B(_3756_), .C(_3794_), .Y(_3795_) );
NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_3__2_), .B(_3730__bF_buf0), .Y(_3796_) );
NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_6__2_), .B(_3706__bF_buf1), .Y(_3797_) );
AOI22X1 AOI22X1_812 ( .gnd(gnd), .vdd(vdd), .A(_3721_), .B(w_mem_inst_w_mem_8__2_), .C(w_mem_inst_w_mem_4__2_), .D(_3740__bF_buf2), .Y(_3798_) );
NAND3X1 NAND3X1_317 ( .gnd(gnd), .vdd(vdd), .A(_3796_), .B(_3797_), .C(_3798_), .Y(_3799_) );
AOI22X1 AOI22X1_813 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_15__2_), .B(_3738__bF_buf1), .C(w_mem_inst_w_mem_7__2_), .D(_3736__bF_buf2), .Y(_3800_) );
NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_2__2_), .B(_3700__bF_buf1), .Y(_3801_) );
NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_11__2_), .B(_3745__bF_buf3), .Y(_3802_) );
NAND3X1 NAND3X1_318 ( .gnd(gnd), .vdd(vdd), .A(_3802_), .B(_3801_), .C(_3800_), .Y(_3803_) );
NOR3X1 NOR3X1_95 ( .gnd(gnd), .vdd(vdd), .A(_3795_), .B(_3803_), .C(_3799_), .Y(_3804_) );
AOI22X1 AOI22X1_814 ( .gnd(gnd), .vdd(vdd), .A(_3692__bF_buf2), .B(_3781_), .C(_3792_), .D(_3804_), .Y(w_2_) );
XNOR2X1 XNOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_8__2_), .B(w_mem_inst_w_mem_13__2_), .Y(_3805_) );
XNOR2X1 XNOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(w_mem_inst_w_mem_0__2_), .B(w_mem_inst_w_mem_2__2_), .Y(_3806_) );
endmodule
